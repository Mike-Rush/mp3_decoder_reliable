// 
//  MAC_MP3: A Low Energy Implementation of an Audio Decoder
//
//  Copyright (C) 2007 McMaster University
// 
//==============================================================================
// 
// This file is part of MAC_MP3
// 
// MAC_MP3 is distributed in the hope that it will be useful for further research,
// but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY
// or FITNESS FOR A PARTICULAR PURPOSE. MAC_MP3 is free; you can redistribute it
// and/or modify it provided that proper reference is provided to the authors. See
// the documents included in the "doc" folder for further details.
//
//==============================================================================


`timescale 1ns / 100ps

`include "defines.v"

module mac_ram(clock, mem_en, address, data_out);

input clock;
input mem_en;
input [`ADDRESS_WIDTH-1:0] address;
output [`DATA_WIDTH-1:0] data_out;

// Instantiate the RAM
RAMB16_S18 instance_mac_ram_RAMB16_S18 (
	.DO(data_out),
	.DOP(),
	.ADDR(address),
	.CLK(clock),
	.DI(16'h0),
	.DIP(2'b00),
	.EN(mem_en),
	.SSR(1'b0),
	.WE(1'b0)
);

// This is frame 1, gr 0, ch 0
// This is randomly generated
// This is sample 9-17
// synthesis attribute INIT_00 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003BAED3AAF94DD38B708078480E65738DF7A5C"
// This is sample 18-26
// synthesis attribute INIT_01 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003C1C466567A451617C84C27BCA82DC9D858A5"
// This is sample 27-35
// synthesis attribute INIT_02 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300036FD8D006D2B25C5587338D3CA232A4443477"
// This is sample 36-44
// synthesis attribute INIT_03 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300038D2FB7F229942FA187AFDAC844B59B27E749"
// This is sample 45-53
// synthesis attribute INIT_04 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003CB7B8E4AE61D5A857E2F6254F44307721D0C"
// This is sample 54-62
// synthesis attribute INIT_05 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003A47176E43EE2A447A2CE0B8E3DB414433727"
// This is sample 63-71
// synthesis attribute INIT_06 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300037CC6A274ED23FB4384C68FA48409E2841820"
// This is sample 72-80
// synthesis attribute INIT_07 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003FBC9C802F9A110D459DEC14FAF8ADFD3D4B9"
// This is sample 81-89
// synthesis attribute INIT_08 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300033F14465BF9353184AE3546CA5786D13669DF"
// This is sample 90-98
// synthesis attribute INIT_09 of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000398EEA4A603D5714760C69ACA99CDF17E4842"
// This is sample 99-107
// synthesis attribute INIT_0A of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003DF3DBF8D15CEE26B062624E0FACE9A344ACF"
// This is sample 108-116
// synthesis attribute INIT_0B of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003C5BEF8DEA8DBE81C902AFF08816087725944"
// This is sample 117-125
// synthesis attribute INIT_0C of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003D31DF376926C8E6C7EC8A438B54497D3673F"
// This is sample 126-134
// synthesis attribute INIT_0D of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003EB403CB229727065173024D18BDCC7F04610"
// This is sample 135-143
// synthesis attribute INIT_0E of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000335C1EE07B45FFB2631FD184C90F26C27DEC5"
// This is sample 144-152
// synthesis attribute INIT_0F of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003A4898A50B6AA620E01BA9E2669081A442C72"
// This is sample 153-161
// synthesis attribute INIT_10 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003918100507B74BD009CFD99F0F05D9C142050"
// This is sample 162-170
// synthesis attribute INIT_11 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300032EFABB8D374D642E02942EF5E86C47ADE1EF"
// This is sample 171-179
// synthesis attribute INIT_12 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003121D82C4A47AB8C1E1AB8C7E0DF5EF373534"
// This is sample 180-188
// synthesis attribute INIT_13 of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000393EAD369327D0D0AFC8E72861FC3E1304845"
// This is sample 189-197
// synthesis attribute INIT_14 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003D41F6E4EF7C8EB3D902E858F40319643EAF1"
// This is sample 198-206
// synthesis attribute INIT_15 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003E59125E96DFD209A9DD9EE472D2D75E1523A"
// This is sample 207-215
// synthesis attribute INIT_16 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003FB1E5E3D22C71E6BBA519408CA8730289F7E"
// This is sample 216-224
// synthesis attribute INIT_17 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003A4EFB6D290BEEFA661E8E6C4B6FE7EFF9348"
// This is sample 225-233
// synthesis attribute INIT_18 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300035AB75E984EAD0F40DA2608402F8932B54B7D"
// This is sample 234-242
// synthesis attribute INIT_19 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300033D3EB68653AD7E881DD81FF97FCBC4B5A749"
// This is sample 243-251
// synthesis attribute INIT_1A of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003A963F8CA421E9173CFB58085DE351D97B71E"
// This is sample 252-260
// synthesis attribute INIT_1B of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300039ABD7DCB036F8732FC81834C7523F60FBA7B"
// This is sample 261-269
// synthesis attribute INIT_1C of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000336D02CDCDCBD2604A08BE61563100569216B"
// This is sample 270-278
// synthesis attribute INIT_1D of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003B4011BDA3380ECA47C652815EFB4261F9E7D"
// This is sample 279-287
// synthesis attribute INIT_1E of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003A3435AAB41E1275C371CD0EC9CA35261B08A"
// This is sample 288-296
// synthesis attribute INIT_1F of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300034E48FE38CEE8C41B9B9E83EAD8735E02B505"
// This is sample 297-305
// synthesis attribute INIT_20 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003537357B9FE3D78CD5B523E651E3DB731691C"
// This is sample 306-314
// synthesis attribute INIT_21 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300037FA10C8B9B3610623993622C71A6D6E9D7A2"
// This is sample 315-323
// synthesis attribute INIT_22 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003E5CCB457F36D80EBEC7E24A1B441B8023CA9"
// This is sample 324-332
// synthesis attribute INIT_23 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003DB3C015AC3D5A30DC52FBBB64D767943C3FE"
// This is sample 333-341
// synthesis attribute INIT_24 of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000335DE9C1571E94F3E053E1E194D8011716929"
// This is sample 342-350
// synthesis attribute INIT_25 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003678B1283B3188BCEB2052D7E4FB58FD6A5AF"
// This is sample 351-359
// synthesis attribute INIT_26 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003BE53FC0961457BB3511685C594469063DED9"
// This is sample 360-368
// synthesis attribute INIT_27 of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000392A82446710D99A65A513E03DDF978504E58"
// This is sample 369-377
// synthesis attribute INIT_28 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300037B900843992B1F2C51F6D8E3149F49CC770E"
// This is sample 378-386
// synthesis attribute INIT_29 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003A655A3CC3C30EAFB19ADBF308473A66E66C7"
// This is sample 387-395
// synthesis attribute INIT_2A of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003B179B4D704A46963DA188A936FA41B5C56D2"
// This is sample 396-404
// synthesis attribute INIT_2B of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003F7B0AA0F797B658E583A909DD0BE040CB689"
// This is sample 405-413
// synthesis attribute INIT_2C of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003274116D5D2F2FFEBA7EE16EB7D346F04842C"
// This is sample 414-422
// synthesis attribute INIT_2D of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300036C90C0230C9748BBC86CE6E5AF6CCA0B5BFB"
// This is sample 423-431
// synthesis attribute INIT_2E of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000365F9AF89E8BCC80D57653023FCBEA1889350"
// This is sample 432-440
// synthesis attribute INIT_2F of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300037F2D93CDBB86BE5C1278FD0B086C87C2CE6D"
// This is sample 441-449
// synthesis attribute INIT_30 of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000373B3A7E895D04F5209913393ECDF0A349679"
// This is sample 450-458
// synthesis attribute INIT_31 of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000349517BF9F9273C6CDBC4603F6BA917862C91"
// This is sample 459-467
// synthesis attribute INIT_32 of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000344E9F6A6073489542A3BA9FD611101F47202"
// This is sample 468-476
// synthesis attribute INIT_33 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300030996477F9B75C2CE451EF6A299AC7E8D5269"
// This is sample 477-485
// synthesis attribute INIT_34 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003F8D017E21EC1701FDC59D3EE451E871C881E"
// This is sample 486-494
// synthesis attribute INIT_35 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003056CD9203B958B86E9924216CE9F15A85C3E"
// This is sample 495-503
// synthesis attribute INIT_36 of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003033E2356DE1819CC8889993DB573926B2798"
// This is sample 504-512
// synthesis attribute INIT_37 of instance_mac_ram_RAMB16_S18 is "256'h000300030003000300030003000371D06762865936CB6A00256A8EA94244E5AE"
// This is sample 513-521
// synthesis attribute INIT_38 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300034B99AD86FE84CCE590B2603AD4FD70223C89"
// This is sample 522-530
// synthesis attribute INIT_39 of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300038A006B3125BC4508937E0BEF18304EE66912"
// This is sample 531-539
// synthesis attribute INIT_3A of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003F2B144FFCEAFAECB48D1E84D34744E014493"
// This is sample 540-548
// synthesis attribute INIT_3B of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300039B0CC4D9AF6349CBA33275140827108A465F"
// This is sample 549-557
// synthesis attribute INIT_3C of instance_mac_ram_RAMB16_S18 is "256'h00030003000300030003000300031196EBBE39608519153181A3E682003A5D7E"
// This is sample 558-566
// synthesis attribute INIT_3D of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003F4A1453AFA1825F8D86A048D6FF071D59015"
// This is sample 567-575
// synthesis attribute INIT_3E of instance_mac_ram_RAMB16_S18 is "256'h0003000300030003000300030003FD19C809E7EA65D21C1043D478DA625F889A"
// This is sample 0-8
// synthesis attribute INIT_3F of instance_mac_ram_RAMB16_S18 is "256'h0000000000000000000000000000DA95CF8FBB74432ADF49191513C1296EA62E"

// synthesis translate_off

defparam instance_mac_ram_RAMB16_S18.INIT_00 = 256'h0003_0003_0003_0003_0003_0003_0003_BAED_3AAF_94DD_38B7_0807_8480_E657_38DF_7A5C;
defparam instance_mac_ram_RAMB16_S18.INIT_01 = 256'h0003_0003_0003_0003_0003_0003_0003_C1C4_6656_7A45_1617_C84C_27BC_A82D_C9D8_58A5;
defparam instance_mac_ram_RAMB16_S18.INIT_02 = 256'h0003_0003_0003_0003_0003_0003_0003_6FD8_D006_D2B2_5C55_8733_8D3C_A232_A444_3477;
defparam instance_mac_ram_RAMB16_S18.INIT_03 = 256'h0003_0003_0003_0003_0003_0003_0003_8D2F_B7F2_2994_2FA1_87AF_DAC8_44B5_9B27_E749;
defparam instance_mac_ram_RAMB16_S18.INIT_04 = 256'h0003_0003_0003_0003_0003_0003_0003_CB7B_8E4A_E61D_5A85_7E2F_6254_F443_0772_1D0C;
defparam instance_mac_ram_RAMB16_S18.INIT_05 = 256'h0003_0003_0003_0003_0003_0003_0003_A471_76E4_3EE2_A447_A2CE_0B8E_3DB4_1443_3727;
defparam instance_mac_ram_RAMB16_S18.INIT_06 = 256'h0003_0003_0003_0003_0003_0003_0003_7CC6_A274_ED23_FB43_84C6_8FA4_8409_E284_1820;
defparam instance_mac_ram_RAMB16_S18.INIT_07 = 256'h0003_0003_0003_0003_0003_0003_0003_FBC9_C802_F9A1_10D4_59DE_C14F_AF8A_DFD3_D4B9;
defparam instance_mac_ram_RAMB16_S18.INIT_08 = 256'h0003_0003_0003_0003_0003_0003_0003_3F14_465B_F935_3184_AE35_46CA_5786_D136_69DF;
defparam instance_mac_ram_RAMB16_S18.INIT_09 = 256'h0003_0003_0003_0003_0003_0003_0003_98EE_A4A6_03D5_7147_60C6_9ACA_99CD_F17E_4842;
defparam instance_mac_ram_RAMB16_S18.INIT_0A = 256'h0003_0003_0003_0003_0003_0003_0003_DF3D_BF8D_15CE_E26B_0626_24E0_FACE_9A34_4ACF;
defparam instance_mac_ram_RAMB16_S18.INIT_0B = 256'h0003_0003_0003_0003_0003_0003_0003_C5BE_F8DE_A8DB_E81C_902A_FF08_8160_8772_5944;
defparam instance_mac_ram_RAMB16_S18.INIT_0C = 256'h0003_0003_0003_0003_0003_0003_0003_D31D_F376_926C_8E6C_7EC8_A438_B544_97D3_673F;
defparam instance_mac_ram_RAMB16_S18.INIT_0D = 256'h0003_0003_0003_0003_0003_0003_0003_EB40_3CB2_2972_7065_1730_24D1_8BDC_C7F0_4610;
defparam instance_mac_ram_RAMB16_S18.INIT_0E = 256'h0003_0003_0003_0003_0003_0003_0003_35C1_EE07_B45F_FB26_31FD_184C_90F2_6C27_DEC5;
defparam instance_mac_ram_RAMB16_S18.INIT_0F = 256'h0003_0003_0003_0003_0003_0003_0003_A489_8A50_B6AA_620E_01BA_9E26_6908_1A44_2C72;
defparam instance_mac_ram_RAMB16_S18.INIT_10 = 256'h0003_0003_0003_0003_0003_0003_0003_9181_0050_7B74_BD00_9CFD_99F0_F05D_9C14_2050;
defparam instance_mac_ram_RAMB16_S18.INIT_11 = 256'h0003_0003_0003_0003_0003_0003_0003_2EFA_BB8D_374D_642E_0294_2EF5_E86C_47AD_E1EF;
defparam instance_mac_ram_RAMB16_S18.INIT_12 = 256'h0003_0003_0003_0003_0003_0003_0003_121D_82C4_A47A_B8C1_E1AB_8C7E_0DF5_EF37_3534;
defparam instance_mac_ram_RAMB16_S18.INIT_13 = 256'h0003_0003_0003_0003_0003_0003_0003_93EA_D369_327D_0D0A_FC8E_7286_1FC3_E130_4845;
defparam instance_mac_ram_RAMB16_S18.INIT_14 = 256'h0003_0003_0003_0003_0003_0003_0003_D41F_6E4E_F7C8_EB3D_902E_858F_4031_9643_EAF1;
defparam instance_mac_ram_RAMB16_S18.INIT_15 = 256'h0003_0003_0003_0003_0003_0003_0003_E591_25E9_6DFD_209A_9DD9_EE47_2D2D_75E1_523A;
defparam instance_mac_ram_RAMB16_S18.INIT_16 = 256'h0003_0003_0003_0003_0003_0003_0003_FB1E_5E3D_22C7_1E6B_BA51_9408_CA87_3028_9F7E;
defparam instance_mac_ram_RAMB16_S18.INIT_17 = 256'h0003_0003_0003_0003_0003_0003_0003_A4EF_B6D2_90BE_EFA6_61E8_E6C4_B6FE_7EFF_9348;
defparam instance_mac_ram_RAMB16_S18.INIT_18 = 256'h0003_0003_0003_0003_0003_0003_0003_5AB7_5E98_4EAD_0F40_DA26_0840_2F89_32B5_4B7D;
defparam instance_mac_ram_RAMB16_S18.INIT_19 = 256'h0003_0003_0003_0003_0003_0003_0003_3D3E_B686_53AD_7E88_1DD8_1FF9_7FCB_C4B5_A749;
defparam instance_mac_ram_RAMB16_S18.INIT_1A = 256'h0003_0003_0003_0003_0003_0003_0003_A963_F8CA_421E_9173_CFB5_8085_DE35_1D97_B71E;
defparam instance_mac_ram_RAMB16_S18.INIT_1B = 256'h0003_0003_0003_0003_0003_0003_0003_9ABD_7DCB_036F_8732_FC81_834C_7523_F60F_BA7B;
defparam instance_mac_ram_RAMB16_S18.INIT_1C = 256'h0003_0003_0003_0003_0003_0003_0003_36D0_2CDC_DCBD_2604_A08B_E615_6310_0569_216B;
defparam instance_mac_ram_RAMB16_S18.INIT_1D = 256'h0003_0003_0003_0003_0003_0003_0003_B401_1BDA_3380_ECA4_7C65_2815_EFB4_261F_9E7D;
defparam instance_mac_ram_RAMB16_S18.INIT_1E = 256'h0003_0003_0003_0003_0003_0003_0003_A343_5AAB_41E1_275C_371C_D0EC_9CA3_5261_B08A;
defparam instance_mac_ram_RAMB16_S18.INIT_1F = 256'h0003_0003_0003_0003_0003_0003_0003_4E48_FE38_CEE8_C41B_9B9E_83EA_D873_5E02_B505;
defparam instance_mac_ram_RAMB16_S18.INIT_20 = 256'h0003_0003_0003_0003_0003_0003_0003_5373_57B9_FE3D_78CD_5B52_3E65_1E3D_B731_691C;
defparam instance_mac_ram_RAMB16_S18.INIT_21 = 256'h0003_0003_0003_0003_0003_0003_0003_7FA1_0C8B_9B36_1062_3993_622C_71A6_D6E9_D7A2;
defparam instance_mac_ram_RAMB16_S18.INIT_22 = 256'h0003_0003_0003_0003_0003_0003_0003_E5CC_B457_F36D_80EB_EC7E_24A1_B441_B802_3CA9;
defparam instance_mac_ram_RAMB16_S18.INIT_23 = 256'h0003_0003_0003_0003_0003_0003_0003_DB3C_015A_C3D5_A30D_C52F_BBB6_4D76_7943_C3FE;
defparam instance_mac_ram_RAMB16_S18.INIT_24 = 256'h0003_0003_0003_0003_0003_0003_0003_35DE_9C15_71E9_4F3E_053E_1E19_4D80_1171_6929;
defparam instance_mac_ram_RAMB16_S18.INIT_25 = 256'h0003_0003_0003_0003_0003_0003_0003_678B_1283_B318_8BCE_B205_2D7E_4FB5_8FD6_A5AF;
defparam instance_mac_ram_RAMB16_S18.INIT_26 = 256'h0003_0003_0003_0003_0003_0003_0003_BE53_FC09_6145_7BB3_5116_85C5_9446_9063_DED9;
defparam instance_mac_ram_RAMB16_S18.INIT_27 = 256'h0003_0003_0003_0003_0003_0003_0003_92A8_2446_710D_99A6_5A51_3E03_DDF9_7850_4E58;
defparam instance_mac_ram_RAMB16_S18.INIT_28 = 256'h0003_0003_0003_0003_0003_0003_0003_7B90_0843_992B_1F2C_51F6_D8E3_149F_49CC_770E;
defparam instance_mac_ram_RAMB16_S18.INIT_29 = 256'h0003_0003_0003_0003_0003_0003_0003_A655_A3CC_3C30_EAFB_19AD_BF30_8473_A66E_66C7;
defparam instance_mac_ram_RAMB16_S18.INIT_2A = 256'h0003_0003_0003_0003_0003_0003_0003_B179_B4D7_04A4_6963_DA18_8A93_6FA4_1B5C_56D2;
defparam instance_mac_ram_RAMB16_S18.INIT_2B = 256'h0003_0003_0003_0003_0003_0003_0003_F7B0_AA0F_797B_658E_583A_909D_D0BE_040C_B689;
defparam instance_mac_ram_RAMB16_S18.INIT_2C = 256'h0003_0003_0003_0003_0003_0003_0003_2741_16D5_D2F2_FFEB_A7EE_16EB_7D34_6F04_842C;
defparam instance_mac_ram_RAMB16_S18.INIT_2D = 256'h0003_0003_0003_0003_0003_0003_0003_6C90_C023_0C97_48BB_C86C_E6E5_AF6C_CA0B_5BFB;
defparam instance_mac_ram_RAMB16_S18.INIT_2E = 256'h0003_0003_0003_0003_0003_0003_0003_65F9_AF89_E8BC_C80D_5765_3023_FCBE_A188_9350;
defparam instance_mac_ram_RAMB16_S18.INIT_2F = 256'h0003_0003_0003_0003_0003_0003_0003_7F2D_93CD_BB86_BE5C_1278_FD0B_086C_87C2_CE6D;
defparam instance_mac_ram_RAMB16_S18.INIT_30 = 256'h0003_0003_0003_0003_0003_0003_0003_73B3_A7E8_95D0_4F52_0991_3393_ECDF_0A34_9679;
defparam instance_mac_ram_RAMB16_S18.INIT_31 = 256'h0003_0003_0003_0003_0003_0003_0003_4951_7BF9_F927_3C6C_DBC4_603F_6BA9_1786_2C91;
defparam instance_mac_ram_RAMB16_S18.INIT_32 = 256'h0003_0003_0003_0003_0003_0003_0003_44E9_F6A6_0734_8954_2A3B_A9FD_6111_01F4_7202;
defparam instance_mac_ram_RAMB16_S18.INIT_33 = 256'h0003_0003_0003_0003_0003_0003_0003_0996_477F_9B75_C2CE_451E_F6A2_99AC_7E8D_5269;
defparam instance_mac_ram_RAMB16_S18.INIT_34 = 256'h0003_0003_0003_0003_0003_0003_0003_F8D0_17E2_1EC1_701F_DC59_D3EE_451E_871C_881E;
defparam instance_mac_ram_RAMB16_S18.INIT_35 = 256'h0003_0003_0003_0003_0003_0003_0003_056C_D920_3B95_8B86_E992_4216_CE9F_15A8_5C3E;
defparam instance_mac_ram_RAMB16_S18.INIT_36 = 256'h0003_0003_0003_0003_0003_0003_0003_033E_2356_DE18_19CC_8889_993D_B573_926B_2798;
defparam instance_mac_ram_RAMB16_S18.INIT_37 = 256'h0003_0003_0003_0003_0003_0003_0003_71D0_6762_8659_36CB_6A00_256A_8EA9_4244_E5AE;
defparam instance_mac_ram_RAMB16_S18.INIT_38 = 256'h0003_0003_0003_0003_0003_0003_0003_4B99_AD86_FE84_CCE5_90B2_603A_D4FD_7022_3C89;
defparam instance_mac_ram_RAMB16_S18.INIT_39 = 256'h0003_0003_0003_0003_0003_0003_0003_8A00_6B31_25BC_4508_937E_0BEF_1830_4EE6_6912;
defparam instance_mac_ram_RAMB16_S18.INIT_3A = 256'h0003_0003_0003_0003_0003_0003_0003_F2B1_44FF_CEAF_AECB_48D1_E84D_3474_4E01_4493;
defparam instance_mac_ram_RAMB16_S18.INIT_3B = 256'h0003_0003_0003_0003_0003_0003_0003_9B0C_C4D9_AF63_49CB_A332_7514_0827_108A_465F;
defparam instance_mac_ram_RAMB16_S18.INIT_3C = 256'h0003_0003_0003_0003_0003_0003_0003_1196_EBBE_3960_8519_1531_81A3_E682_003A_5D7E;
defparam instance_mac_ram_RAMB16_S18.INIT_3D = 256'h0003_0003_0003_0003_0003_0003_0003_F4A1_453A_FA18_25F8_D86A_048D_6FF0_71D5_9015;
defparam instance_mac_ram_RAMB16_S18.INIT_3E = 256'h0003_0003_0003_0003_0003_0003_0003_FD19_C809_E7EA_65D2_1C10_43D4_78DA_625F_889A;
defparam instance_mac_ram_RAMB16_S18.INIT_3F = 256'h0000_0000_0000_0000_0000_0000_0000_DA95_CF8F_BB74_432A_DF49_1915_13C1_296E_A62E;

// synthesis translate_on


endmodule
