// 
//  MAC_MP3: A Low Energy Implementation of an Audio Decoder
//
//  Copyright (C) 2007 McMaster University
// 
//==============================================================================
// 
// This file is part of MAC_MP3
// 
// MAC_MP3 is distributed in the hope that it will be useful for further research,
// but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY
// or FITNESS FOR A PARTICULAR PURPOSE. MAC_MP3 is free; you can redistribute it
// and/or modify it provided that proper reference is provided to the authors. See
// the documents included in the "doc" folder for further details.
//
//==============================================================================


`timescale 1ns / 100ps

`include "../defines.v"

module polyphase_sample_buffer(clock, mem_en, wr_en, address, data_in ,data_out);

input clock;
input mem_en;
input wr_en;
input [`ADDRESS_WIDTH-1:0] address;
input [`DATA_WIDTH-1:0] data_in;
output [`DATA_WIDTH-1:0] data_out;

// Instantiate the RAM
RAMB16_S18 instance_polyphase_sample_buffer_RAMB16_S18(
	.DO(data_out),
	.DOP(),
	.ADDR(address),
	.CLK(clock),
	.DI(data_in),
	.DIP(2'b00),
	.EN(mem_en),
	.SSR(1'b0),
	.WE(wr_en)
);

// synthesis attribute INIT_00 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_01 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_02 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_03 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_04 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_05 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_06 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_07 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_08 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_09 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0A of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0B of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0C of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0D of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0E of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0F of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_10 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_11 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_12 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_13 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_14 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_15 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_16 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_17 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_18 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_19 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1A of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1B of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1C of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1D of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1E of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1F of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_20 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_21 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_22 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_23 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_24 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_25 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_26 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_27 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_28 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_29 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2A of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2B of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2C of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2D of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2E of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2F of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_30 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_31 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_32 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_33 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_34 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_35 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_36 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_37 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_38 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_39 of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3A of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3B of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3C of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3D of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3E of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3F of instance_polyphase_sample_buffer_RAMB16_S18 is "256'h0000000000000000000000000000000000000000000000000000000000000000"

// synthesis translate_off

defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_polyphase_sample_buffer_RAMB16_S18.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// synthesis translate_on


endmodule
