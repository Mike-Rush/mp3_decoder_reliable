// 
//  MAC_MP3: A Low Energy Implementation of an Audio Decoder
//
//  Copyright (C) 2007 McMaster University
// 
//==============================================================================
// 
// This file is part of MAC_MP3
// 
// MAC_MP3 is distributed in the hope that it will be useful for further research,
// but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY
// or FITNESS FOR A PARTICULAR PURPOSE. MAC_MP3 is free; you can redistribute it
// and/or modify it provided that proper reference is provided to the authors. See
// the documents included in the "doc" folder for further details.
//
//==============================================================================



`timescale 1 ns / 100 ps

`include "defines.v"

module antialias_imdct_coefficient (
	clock,
	CH0_mem_en,
	CH0_address,
	CH0_data_out,
	CH1_mem_en,
	CH1_address,
	CH1_data_out
);

input clock;
input CH0_mem_en, CH1_mem_en;
input [`ADDRESS_WIDTH-1:0] CH0_address, CH1_address;
output [`DATA_WIDTH-1:0] CH0_data_out, CH1_data_out;

// Instantiate the RAM



	RAMB16_S18_S18 antialias_imdct_coefficient_RAM (
    .DOA(CH0_data_out),
    .DOPA(),
    .ADDRA(CH0_address),
    .CLKA(clock),
    .DIA(16'h0000),
    .DIPA(2'b00),
    .ENA(CH0_mem_en),
    .SSRA(1'b0),
    .WEA(1'b0),

	 

	 .DOB(CH1_data_out),
    .DOPB(),

    .ADDRB(CH1_address),
    .CLKB(clock),
    .DIB(16'h0000),
    .DIPB(2'b00),
    .ENB(CH1_mem_en),
    .SSRB(1'b0),
	 .WEB(1'b0)
  );


// COS coefficient for IMDCT for normal block (0-647)...
// Coe i = 0, k = 0-17
// synthesis attribute INIT_00 of antialias_imdct_coefficient_RAM is "256'h35FA1D8DC4DFECC13E7B085AC00F02CA3F73F225C2F6187D38C4DD9CCD392B3C"
// Coe i = 18, k = 0-17
// synthesis attribute INIT_01 of antialias_imdct_coefficient_RAM is "256'hE782C2F60DDA3F73FD35C00FF7A53E7B133EC4DFE27235FA26F5D0D0D0D0D90A"
// Coe i = 1, k = 0-17
// synthesis attribute INIT_02 of antialias_imdct_coefficient_RAM is "256'hD90A3B20085AC08C187D32C6CD39E7823F73F7A5C4DF26F5D4C3CD39226338C4"
// Coe i = 19, k = 0-17
// synthesis attribute INIT_03 of antialias_imdct_coefficient_RAM is "256'hC08CF7A53B2026F5D90AC4DF085A3F73187DCD3932C6187DC08C085A3B20D90A"
// Coe i = 2, k = 0-17
// synthesis attribute INIT_04 of antialias_imdct_coefficient_RAM is "256'hCD3938C402CAC4DF2F2F133EC08C226326F63B20F7A5C08CE78232C632C6E782"
// Coe i = 20, k = 0-17
// synthesis attribute INIT_05 of antialias_imdct_coefficient_RAM is "256'hC00FE7822B3C3D09085ACA05CA05F7A53D09D4C3E7823FF0E272D90A3E7BF225"
// Coe i = 3, k = 0-17
// synthesis attribute INIT_06 of antialias_imdct_coefficient_RAM is "256'h0DDA2B3CC08C1D8DDD9CC08CECC12F2F3B2002CAC73BCD390DDA3E7B26F5E272"
// Coe i = 21, k = 0-17
// synthesis attribute INIT_07 of antialias_imdct_coefficient_RAM is "256'hF7A5C73B38C4F7A5D0D03E7BE782DD9C3FF0D90AECC13D09CD39FD3535FAC4DF"
// synthesis attribute INIT_08 of antialias_imdct_coefficient_RAM is "256'h1D8D3F732B3CF225C4DFCA05FD3532C63D09133ED90AC00FDD9C187D3E7B2F2F"
// Coe i = 4, k = 0-17
// synthesis attribute INIT_09 of antialias_imdct_coefficient_RAM is "256'h187DC4DF3B20E782E7823B20C4DF187D187DC4DF3B20E782E7823B20C4DF187D"
// Coe i = 22, k = 0-17
// synthesis attribute INIT_0A of antialias_imdct_coefficient_RAM is "256'h187D3B203B20187DE782C4DFC4DFE782187D3B203B20187DE782C4DFC4DF187D"
// Coe i = 5, k = 0-17
// synthesis attribute INIT_0B of antialias_imdct_coefficient_RAM is "256'hD4C3085A1D8DC73B3F73D0D00DDA187DCA053FF0CD39133EE782C4DFC4DFE782"
// Coe i = 23, k = 0-17
// synthesis attribute INIT_0C of antialias_imdct_coefficient_RAM is "256'hC73BE272085A2B3C3E7B3B202263FD35D90AC2F63D09D90A02CA2263C4DF3E7B"
// Coe i = 6, k = 0-17
// synthesis attribute INIT_0D of antialias_imdct_coefficient_RAM is "256'h085A133ED4C33B20C00F38C4D90A0DDA133E32C63FF035FA187DF225D0D0C08C"
// Coe i = 24, k = 0-17
// synthesis attribute INIT_0E of antialias_imdct_coefficient_RAM is "256'h2F2F187DFD35E272CD39C184C18432C6E27202CA187DD0D03D09C08C35FADD9C"
// Coe i = 7, k = 0-17
// synthesis attribute INIT_0F of antialias_imdct_coefficient_RAM is "256'hCD3926F5E782085AF225D90AC73BC00FC4DFD4C3ECC1085A226335FA3F733D09"
// Coe i = 25, k = 0-17
// synthesis attribute INIT_10 of antialias_imdct_coefficient_RAM is "256'hC4DFC08C3F73C4DF32C6D90A187DF7A5F7A5187DD90A32C6C4DF3F73C08C3B20"
// synthesis attribute INIT_11 of antialias_imdct_coefficient_RAM is "256'h085A187D26F532C63B203F733F733B2032C626F5187D085AF7A5E782D90ACD39"
// Coe i = 8, k = 0-17
// synthesis attribute INIT_12 of antialias_imdct_coefficient_RAM is "256'hC1843D09C4DF38C4CA0532C6D0D02B3CD90A2263E272187DECC10DDAF7A502CA"
// Coe i = 26, k = 0-17
// synthesis attribute INIT_13 of antialias_imdct_coefficient_RAM is "256'hE782E272DD9CD90AD4C3D0D0CD39CA05C73BC4DFC2F6C184C08CC00FC00F3F73"
// Coe i = 9, k = 0-17
// synthesis attribute INIT_14 of antialias_imdct_coefficient_RAM is "256'h35FACD392F2FD4C326F5DD9C1D8DE782133EF225085AFD35FD35F7A5F225ECC1"
// Coe i = 27, k = 0-17
// synthesis attribute INIT_15 of antialias_imdct_coefficient_RAM is "256'hD4C3D0D0CD39CA05C73BC4DFC2F6C184C08CC00F3FF0C08C3E7BC2F63B20C73B"
// Coe i = 10, k = 0-17
// synthesis attribute INIT_16 of antialias_imdct_coefficient_RAM is "256'h3B20C08C3F73C4DF32C6D90A187DF7A5FD35F7A5F225ECC1E782E272DD9CD90A"
// Coe i = 28, k = 0-17
// synthesis attribute INIT_17 of antialias_imdct_coefficient_RAM is "256'hF7A5E782D90ACD39C4DFC08CC08C3B20CD3926F5E782085A085AE78226F5CD39"
// Coe i = 11, k = 0-17
// synthesis attribute INIT_18 of antialias_imdct_coefficient_RAM is "256'h3FF0C73B26F5F225085A187D26F532C63B203F733F733B2032C626F5187D085A"
// Coe i = 29, k = 0-17
// synthesis attribute INIT_19 of antialias_imdct_coefficient_RAM is "256'hCD39C1843E7BCD391D8DFD35E7822F2FC2F63F73CA052263F7A5ECC12B3CC4DF"
// synthesis attribute INIT_1A of antialias_imdct_coefficient_RAM is "256'hF225D90AC73BC00FC4DFD4C3ECC1085A226335FA3F733D092F2F187DFD35E272"
// Coe i = 12, k = 0-17
// synthesis attribute INIT_1B of antialias_imdct_coefficient_RAM is "256'hFD35DD9C3B20C1842B3CF7A5E27238C4C08C2F2FF225E78235FAC00F32C6ECC1"
// Coe i = 30, k = 0-17
// synthesis attribute INIT_1C of antialias_imdct_coefficient_RAM is "256'h187DF225D0D0C08CC73BE272085A2B3C3E7B3B202263FD35D90AC2F6C2F626F5"
// Coe i = 13, k = 0-17
// synthesis attribute INIT_1D of antialias_imdct_coefficient_RAM is "256'h187DC4DF3B20E782E7823B20C4DF187D187DC4DF3B20E782133E32C63FF035FA"
// Coe i = 31, k = 0-17
// synthesis attribute INIT_1E of antialias_imdct_coefficient_RAM is "256'hE782C4DFC4DFE782187D3B203B20187DE782C4DF3B20E782E7823B20C4DF187D"
// Coe i = 14, k = 0-17
// synthesis attribute INIT_1F of antialias_imdct_coefficient_RAM is "256'h32C602CACA053B20F225D4C33F73E272E782C4DFC4DFE782187D3B203B20187D"
// Coe i = 32, k = 0-17
// synthesis attribute INIT_20 of antialias_imdct_coefficient_RAM is "256'hDD9C187D3E7B2F2FF7A5C73BC73B085A2F2FC184187D2263C00F26F5133EC2F6"
// Coe i = 15, k = 0-17
// synthesis attribute INIT_21 of antialias_imdct_coefficient_RAM is "256'hD0D0ECC13F73DD9C1D8D3F732B3CF225C4DFCA05FD3532C63D09133ED90AC00F"
// Coe i = 33, k = 0-17
// synthesis attribute INIT_22 of antialias_imdct_coefficient_RAM is "256'h085ACA0535FA085AC2F62B3C187DC00F1D8D26F5C1840DDA32C6C73BFD353B20"
// synthesis attribute INIT_23 of antialias_imdct_coefficient_RAM is "256'hDD9CC08CECC12F2F3B2002CAC73BCD390DDA3E7B26F5E272C00FE7822B3C3D09"
// Coe i = 16, k = 0-17
// synthesis attribute INIT_24 of antialias_imdct_coefficient_RAM is "256'h3F73F7A5C4DF26F526F5C4DFF7A53F73E782CD3932C6187DC08C085A3B20D90A"
// Coe i = 34, k = 0-17
// synthesis attribute INIT_25 of antialias_imdct_coefficient_RAM is "256'hE78232C632C6E782C08CF7A53B2026F5D90AC4DF085A3F73187DCD39CD39E782"
// Coe i = 17, k = 0-17
// synthesis attribute INIT_26 of antialias_imdct_coefficient_RAM is "256'hC184F7A53FF0FD35C08C0DDA3D09E782C73B226332C6D4C326F53B20F7A5C08C"
// Coe i = 35, k = 0-17
// synthesis attribute INIT_27 of antialias_imdct_coefficient_RAM is "256'hFD35C00FF7A53E7B133EC4DFE27235FA26F5D0D02F2F26F5CA05E2723B20133E"
// Constant 0 (648-655)...
// synthesis attribute INIT_28 of antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000D4C3CD39226338C4E782C2F60DDA3F73"
// window coefficient for IMDCT block type 2 (656-667)...
// Constant 1 (668-703)...
// synthesis attribute INIT_29 of antialias_imdct_coefficient_RAM is "256'h4000400040004000085A187D26F532C63B203F733F733B2032C626F5187D085A"
// synthesis attribute INIT_2A of antialias_imdct_coefficient_RAM is "256'h4000400040004000400040004000400040004000400040004000400040004000"
// synthesis attribute INIT_2B of antialias_imdct_coefficient_RAM is "256'h4000400040004000400040004000400040004000400040004000400040004000"
// window coefficient for IMDCT block type 0 (704-767)...(index: 0, 18, 1, 19, 2, 20....)
// synthesis attribute INIT_2C of antialias_imdct_coefficient_RAM is "256'h32C626F535FA226338C41D8D3B20187D3D09133E3E7B0DDA3F73085A3FF002CA"
// synthesis attribute INIT_2D of antialias_imdct_coefficient_RAM is "256'h0DDA3E7B133E3D09187D3B201D8D38C4226335FA26F532C62B3C2F2F2F2F2B3C"
// Constant 0 (648-655)...
// synthesis attribute INIT_2E of antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000000000000000000002CA3FF0085A3F73"
// synthesis attribute INIT_2F of antialias_imdct_coefficient_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// window coefficient for IMDCT block type 1 (768-831)...(index: 0, 18, 1, 19, 2, 20....)
// synthesis attribute INIT_30 of antialias_imdct_coefficient_RAM is "256'h3B2026F53F73226340001D8D4000187D4000133E40000DDA4000085A400002CA"
// synthesis attribute INIT_31 of antialias_imdct_coefficient_RAM is "256'h00003E7B00003D0900003B20000038C4085A35FA187D32C626F52F2F32C62B3C"
// Constant 0 (648-655)...
// synthesis attribute INIT_32 of antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000000000000000000000003FF000003F73"
// synthesis attribute INIT_33 of antialias_imdct_coefficient_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// window coefficient for IMDCT block type 3 (832-895)...(index: 0, 18, 1, 19, 2, 20....)
// synthesis attribute INIT_34 of antialias_imdct_coefficient_RAM is "256'h32C6187D35FA085A38C400003B2000003D0900003E7B00003F7300003FF00000"
// synthesis attribute INIT_35 of antialias_imdct_coefficient_RAM is "256'h0DDA4000133E4000187D40001D8D400022633F7326F53B202B3C32C62F2F26F5"
// Constant 0 (648-655)...
// synthesis attribute INIT_36 of antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000000000000000000002CA4000085A4000"
// synthesis attribute INIT_37 of antialias_imdct_coefficient_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// COS coefficient for for IMDCT short block (896-967)...
// synthesis attribute INIT_38 of antialias_imdct_coefficient_RAM is "256'hCD3926F5E782085A3B20E782E7823B20C4DF187DCD39E7823F73F7A5C4DF26F5"
// synthesis attribute INIT_39 of antialias_imdct_coefficient_RAM is "256'h3B20D90AC4DF187D187DC4DF3B20E7823F73C4DF32C6D90A187DF7A5C08C3B20"
// synthesis attribute INIT_3A of antialias_imdct_coefficient_RAM is "256'h187D3B203B20187DE782C4DFD90AC4DF085A3F73187DCD3932C6187DC08C085A"
// synthesis attribute INIT_3B of antialias_imdct_coefficient_RAM is "256'h3B20187DE782C4DFF7A5E782D90ACD39C4DFC08CF7A5E782D90ACD39C4DFC08C"
// Constant -1 (968-999)...
// synthesis attribute INIT_3C of antialias_imdct_coefficient_RAM is "256'hC000C000C000C000C000C000C000C000D90AC4DF085A3F73187DCD39187D3B20"
// synthesis attribute INIT_3D of antialias_imdct_coefficient_RAM is "256'hC000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000"
// CS coefficient (1000-1007)...
// synthesis attribute INIT_3E of antialias_imdct_coefficient_RAM is "256'h3FFF3FFE3FF23FB63EEE3CC6386E36E1C000C000C000C000C000C000C000C000"
// CA coefficient (1008-1015)...
// -CA coefficient (1016-1023)...
// synthesis attribute INIT_3F of antialias_imdct_coefficient_RAM is "256'h003C00E8029F060D0BA4140E1E3020EDFFC3FF17FD60F9F2F45BEBF1E1CFDF12"

// synthesis translate_off

defparam antialias_imdct_coefficient_RAM.INIT_00 = 256'h35FA_1D8D_C4DF_ECC1_3E7B_085A_C00F_02CA_3F73_F225_C2F6_187D_38C4_DD9C_CD39_2B3C;
defparam antialias_imdct_coefficient_RAM.INIT_01 = 256'hE782_C2F6_0DDA_3F73_FD35_C00F_F7A5_3E7B_133E_C4DF_E272_35FA_26F5_D0D0_D0D0_D90A;
defparam antialias_imdct_coefficient_RAM.INIT_02 = 256'hD90A_3B20_085A_C08C_187D_32C6_CD39_E782_3F73_F7A5_C4DF_26F5_D4C3_CD39_2263_38C4;
defparam antialias_imdct_coefficient_RAM.INIT_03 = 256'hC08C_F7A5_3B20_26F5_D90A_C4DF_085A_3F73_187D_CD39_32C6_187D_C08C_085A_3B20_D90A;
defparam antialias_imdct_coefficient_RAM.INIT_04 = 256'hCD39_38C4_02CA_C4DF_2F2F_133E_C08C_2263_26F6_3B20_F7A5_C08C_E782_32C6_32C6_E782;
defparam antialias_imdct_coefficient_RAM.INIT_05 = 256'hC00F_E782_2B3C_3D09_085A_CA05_CA05_F7A5_3D09_D4C3_E782_3FF0_E272_D90A_3E7B_F225;
defparam antialias_imdct_coefficient_RAM.INIT_06 = 256'h0DDA_2B3C_C08C_1D8D_DD9C_C08C_ECC1_2F2F_3B20_02CA_C73B_CD39_0DDA_3E7B_26F5_E272;
defparam antialias_imdct_coefficient_RAM.INIT_07 = 256'hF7A5_C73B_38C4_F7A5_D0D0_3E7B_E782_DD9C_3FF0_D90A_ECC1_3D09_CD39_FD35_35FA_C4DF;
defparam antialias_imdct_coefficient_RAM.INIT_08 = 256'h1D8D_3F73_2B3C_F225_C4DF_CA05_FD35_32C6_3D09_133E_D90A_C00F_DD9C_187D_3E7B_2F2F;
defparam antialias_imdct_coefficient_RAM.INIT_09 = 256'h187D_C4DF_3B20_E782_E782_3B20_C4DF_187D_187D_C4DF_3B20_E782_E782_3B20_C4DF_187D;
defparam antialias_imdct_coefficient_RAM.INIT_0A = 256'h187D_3B20_3B20_187D_E782_C4DF_C4DF_E782_187D_3B20_3B20_187D_E782_C4DF_C4DF_187D;
defparam antialias_imdct_coefficient_RAM.INIT_0B = 256'hD4C3_085A_1D8D_C73B_3F73_D0D0_0DDA_187D_CA05_3FF0_CD39_133E_E782_C4DF_C4DF_E782;
defparam antialias_imdct_coefficient_RAM.INIT_0C = 256'hC73B_E272_085A_2B3C_3E7B_3B20_2263_FD35_D90A_C2F6_3D09_D90A_02CA_2263_C4DF_3E7B;
defparam antialias_imdct_coefficient_RAM.INIT_0D = 256'h085A_133E_D4C3_3B20_C00F_38C4_D90A_0DDA_133E_32C6_3FF0_35FA_187D_F225_D0D0_C08C;
defparam antialias_imdct_coefficient_RAM.INIT_0E = 256'h2F2F_187D_FD35_E272_CD39_C184_C184_32C6_E272_02CA_187D_D0D0_3D09_C08C_35FA_DD9C;
defparam antialias_imdct_coefficient_RAM.INIT_0F = 256'hCD39_26F5_E782_085A_F225_D90A_C73B_C00F_C4DF_D4C3_ECC1_085A_2263_35FA_3F73_3D09;
defparam antialias_imdct_coefficient_RAM.INIT_10 = 256'hC4DF_C08C_3F73_C4DF_32C6_D90A_187D_F7A5_F7A5_187D_D90A_32C6_C4DF_3F73_C08C_3B20;
defparam antialias_imdct_coefficient_RAM.INIT_11 = 256'h085A_187D_26F5_32C6_3B20_3F73_3F73_3B20_32C6_26F5_187D_085A_F7A5_E782_D90A_CD39;
defparam antialias_imdct_coefficient_RAM.INIT_12 = 256'hC184_3D09_C4DF_38C4_CA05_32C6_D0D0_2B3C_D90A_2263_E272_187D_ECC1_0DDA_F7A5_02CA;
defparam antialias_imdct_coefficient_RAM.INIT_13 = 256'hE782_E272_DD9C_D90A_D4C3_D0D0_CD39_CA05_C73B_C4DF_C2F6_C184_C08C_C00F_C00F_3F73;
defparam antialias_imdct_coefficient_RAM.INIT_14 = 256'h35FA_CD39_2F2F_D4C3_26F5_DD9C_1D8D_E782_133E_F225_085A_FD35_FD35_F7A5_F225_ECC1;
defparam antialias_imdct_coefficient_RAM.INIT_15 = 256'hD4C3_D0D0_CD39_CA05_C73B_C4DF_C2F6_C184_C08C_C00F_3FF0_C08C_3E7B_C2F6_3B20_C73B;
defparam antialias_imdct_coefficient_RAM.INIT_16 = 256'h3B20_C08C_3F73_C4DF_32C6_D90A_187D_F7A5_FD35_F7A5_F225_ECC1_E782_E272_DD9C_D90A;
defparam antialias_imdct_coefficient_RAM.INIT_17 = 256'hF7A5_E782_D90A_CD39_C4DF_C08C_C08C_3B20_CD39_26F5_E782_085A_085A_E782_26F5_CD39;
defparam antialias_imdct_coefficient_RAM.INIT_18 = 256'h3FF0_C73B_26F5_F225_085A_187D_26F5_32C6_3B20_3F73_3F73_3B20_32C6_26F5_187D_085A;
defparam antialias_imdct_coefficient_RAM.INIT_19 = 256'hCD39_C184_3E7B_CD39_1D8D_FD35_E782_2F2F_C2F6_3F73_CA05_2263_F7A5_ECC1_2B3C_C4DF;
defparam antialias_imdct_coefficient_RAM.INIT_1A = 256'hF225_D90A_C73B_C00F_C4DF_D4C3_ECC1_085A_2263_35FA_3F73_3D09_2F2F_187D_FD35_E272;
defparam antialias_imdct_coefficient_RAM.INIT_1B = 256'hFD35_DD9C_3B20_C184_2B3C_F7A5_E272_38C4_C08C_2F2F_F225_E782_35FA_C00F_32C6_ECC1;
defparam antialias_imdct_coefficient_RAM.INIT_1C = 256'h187D_F225_D0D0_C08C_C73B_E272_085A_2B3C_3E7B_3B20_2263_FD35_D90A_C2F6_C2F6_26F5;
defparam antialias_imdct_coefficient_RAM.INIT_1D = 256'h187D_C4DF_3B20_E782_E782_3B20_C4DF_187D_187D_C4DF_3B20_E782_133E_32C6_3FF0_35FA;
defparam antialias_imdct_coefficient_RAM.INIT_1E = 256'hE782_C4DF_C4DF_E782_187D_3B20_3B20_187D_E782_C4DF_3B20_E782_E782_3B20_C4DF_187D;
defparam antialias_imdct_coefficient_RAM.INIT_1F = 256'h32C6_02CA_CA05_3B20_F225_D4C3_3F73_E272_E782_C4DF_C4DF_E782_187D_3B20_3B20_187D;
defparam antialias_imdct_coefficient_RAM.INIT_20 = 256'hDD9C_187D_3E7B_2F2F_F7A5_C73B_C73B_085A_2F2F_C184_187D_2263_C00F_26F5_133E_C2F6;
defparam antialias_imdct_coefficient_RAM.INIT_21 = 256'hD0D0_ECC1_3F73_DD9C_1D8D_3F73_2B3C_F225_C4DF_CA05_FD35_32C6_3D09_133E_D90A_C00F;
defparam antialias_imdct_coefficient_RAM.INIT_22 = 256'h085A_CA05_35FA_085A_C2F6_2B3C_187D_C00F_1D8D_26F5_C184_0DDA_32C6_C73B_FD35_3B20;
defparam antialias_imdct_coefficient_RAM.INIT_23 = 256'hDD9C_C08C_ECC1_2F2F_3B20_02CA_C73B_CD39_0DDA_3E7B_26F5_E272_C00F_E782_2B3C_3D09;
defparam antialias_imdct_coefficient_RAM.INIT_24 = 256'h3F73_F7A5_C4DF_26F5_26F5_C4DF_F7A5_3F73_E782_CD39_32C6_187D_C08C_085A_3B20_D90A;
defparam antialias_imdct_coefficient_RAM.INIT_25 = 256'hE782_32C6_32C6_E782_C08C_F7A5_3B20_26F5_D90A_C4DF_085A_3F73_187D_CD39_CD39_E782;
defparam antialias_imdct_coefficient_RAM.INIT_26 = 256'hC184_F7A5_3FF0_FD35_C08C_0DDA_3D09_E782_C73B_2263_32C6_D4C3_26F5_3B20_F7A5_C08C;
defparam antialias_imdct_coefficient_RAM.INIT_27 = 256'hFD35_C00F_F7A5_3E7B_133E_C4DF_E272_35FA_26F5_D0D0_2F2F_26F5_CA05_E272_3B20_133E;
defparam antialias_imdct_coefficient_RAM.INIT_28 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_D4C3_CD39_2263_38C4_E782_C2F6_0DDA_3F73;
defparam antialias_imdct_coefficient_RAM.INIT_29 = 256'h4000_4000_4000_4000_085A_187D_26F5_32C6_3B20_3F73_3F73_3B20_32C6_26F5_187D_085A;
defparam antialias_imdct_coefficient_RAM.INIT_2A = 256'h4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000;
defparam antialias_imdct_coefficient_RAM.INIT_2B = 256'h4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000;
defparam antialias_imdct_coefficient_RAM.INIT_2C = 256'h32C6_26F5_35FA_2263_38C4_1D8D_3B20_187D_3D09_133E_3E7B_0DDA_3F73_085A_3FF0_02CA;
defparam antialias_imdct_coefficient_RAM.INIT_2D = 256'h0DDA_3E7B_133E_3D09_187D_3B20_1D8D_38C4_2263_35FA_26F5_32C6_2B3C_2F2F_2F2F_2B3C;
defparam antialias_imdct_coefficient_RAM.INIT_2E = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_02CA_3FF0_085A_3F73;
defparam antialias_imdct_coefficient_RAM.INIT_2F = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
defparam antialias_imdct_coefficient_RAM.INIT_30 = 256'h3B20_26F5_3F73_2263_4000_1D8D_4000_187D_4000_133E_4000_0DDA_4000_085A_4000_02CA;
defparam antialias_imdct_coefficient_RAM.INIT_31 = 256'h0000_3E7B_0000_3D09_0000_3B20_0000_38C4_085A_35FA_187D_32C6_26F5_2F2F_32C6_2B3C;
defparam antialias_imdct_coefficient_RAM.INIT_32 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_3FF0_0000_3F73;
defparam antialias_imdct_coefficient_RAM.INIT_33 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
defparam antialias_imdct_coefficient_RAM.INIT_34 = 256'h32C6_187D_35FA_085A_38C4_0000_3B20_0000_3D09_0000_3E7B_0000_3F73_0000_3FF0_0000;
defparam antialias_imdct_coefficient_RAM.INIT_35 = 256'h0DDA_4000_133E_4000_187D_4000_1D8D_4000_2263_3F73_26F5_3B20_2B3C_32C6_2F2F_26F5;
defparam antialias_imdct_coefficient_RAM.INIT_36 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_02CA_4000_085A_4000;
defparam antialias_imdct_coefficient_RAM.INIT_37 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
defparam antialias_imdct_coefficient_RAM.INIT_38 = 256'hCD39_26F5_E782_085A_3B20_E782_E782_3B20_C4DF_187D_CD39_E782_3F73_F7A5_C4DF_26F5;
defparam antialias_imdct_coefficient_RAM.INIT_39 = 256'h3B20_D90A_C4DF_187D_187D_C4DF_3B20_E782_3F73_C4DF_32C6_D90A_187D_F7A5_C08C_3B20;
defparam antialias_imdct_coefficient_RAM.INIT_3A = 256'h187D_3B20_3B20_187D_E782_C4DF_D90A_C4DF_085A_3F73_187D_CD39_32C6_187D_C08C_085A;
defparam antialias_imdct_coefficient_RAM.INIT_3B = 256'h3B20_187D_E782_C4DF_F7A5_E782_D90A_CD39_C4DF_C08C_F7A5_E782_D90A_CD39_C4DF_C08C;
defparam antialias_imdct_coefficient_RAM.INIT_3C = 256'hC000_C000_C000_C000_C000_C000_C000_C000_D90A_C4DF_085A_3F73_187D_CD39_187D_3B20;
defparam antialias_imdct_coefficient_RAM.INIT_3D = 256'hC000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000;
defparam antialias_imdct_coefficient_RAM.INIT_3E = 256'h3FFF_3FFE_3FF2_3FB6_3EEE_3CC6_386E_36E1_C000_C000_C000_C000_C000_C000_C000_C000;
defparam antialias_imdct_coefficient_RAM.INIT_3F = 256'h003C_00E8_029F_060D_0BA4_140E_1E30_20ED_FFC3_FF17_FD60_F9F2_F45B_EBF1_E1CF_DF12;

// synthesis translate_on


/*
RAMB16_S18 CH0_antialias_imdct_coefficient_RAM (
	.DO(CH0_data_out),
	.DOP(),
	.ADDR(CH0_address),
	.CLK(clock),
	.DI(16'h0),
	.DIP(2'b00),
	.EN(CH0_mem_en),
	.SSR(1'b0),
	.WE(1'b0)
);

// COS coefficient for IMDCT for normal block (0-647)...
// Coe i = 0, k = 0-17
// synthesis attribute INIT_00 of CH0_antialias_imdct_coefficient_RAM is "256'h35FA1D8DC4DFECC13E7B085AC00F02CA3F73F225C2F6187D38C4DD9CCD392B3C"
// Coe i = 18, k = 0-17
// synthesis attribute INIT_01 of CH0_antialias_imdct_coefficient_RAM is "256'hE782C2F60DDA3F73FD35C00FF7A53E7B133EC4DFE27235FA26F5D0D0D0D0D90A"
// Coe i = 1, k = 0-17
// synthesis attribute INIT_02 of CH0_antialias_imdct_coefficient_RAM is "256'hD90A3B20085AC08C187D32C6CD39E7823F73F7A5C4DF26F5D4C3CD39226338C4"
// Coe i = 19, k = 0-17
// synthesis attribute INIT_03 of CH0_antialias_imdct_coefficient_RAM is "256'hC08CF7A53B2026F5D90AC4DF085A3F73187DCD3932C6187DC08C085A3B20D90A"
// Coe i = 2, k = 0-17
// synthesis attribute INIT_04 of CH0_antialias_imdct_coefficient_RAM is "256'hCD3938C402CAC4DF2F2F133EC08C226326F53B20F7A5C08CE78232C632C6E782"
// Coe i = 20, k = 0-17
// synthesis attribute INIT_05 of CH0_antialias_imdct_coefficient_RAM is "256'hC00FE7822B3C3D09085ACA05CA05F7A53D09D4C3E7823FF0E272D90A3E7BF225"
// Coe i = 3, k = 0-17
// synthesis attribute INIT_06 of CH0_antialias_imdct_coefficient_RAM is "256'h0DDA2B3CC08C1D8DDD9CC08CECC12F2F3B2002CAC73BCD390DDA3E7B26F5E272"
// Coe i = 21, k = 0-17
// synthesis attribute INIT_07 of CH0_antialias_imdct_coefficient_RAM is "256'hF7A5C73B38C4F7A5D0D03E7BE782DD9C3FF0D90AECC13D09CD39FD3535FAC4DF"
// synthesis attribute INIT_08 of CH0_antialias_imdct_coefficient_RAM is "256'h1D8D3F732B3CF225C4DFCA05FD3532C63D09133ED90AC00FDD9C187D3E7B2F2F"
// Coe i = 4, k = 0-17
// synthesis attribute INIT_09 of CH0_antialias_imdct_coefficient_RAM is "256'h187DC4DF3B20E782E7823B20C4DF187D187DC4DF3B20E782E7823B20C4DF187D"
// Coe i = 22, k = 0-17
// synthesis attribute INIT_0A of CH0_antialias_imdct_coefficient_RAM is "256'h187D3B203B20187DE782C4DFC4DFE782187D3B203B20187DE782C4DFC4DF187D"
// Coe i = 5, k = 0-17
// synthesis attribute INIT_0B of CH0_antialias_imdct_coefficient_RAM is "256'hD4C3085A1D8DC73B3F73D0D00DDA187DCA053FF0CD39133EE782C4DFC4DFE782"
// Coe i = 23, k = 0-17
// synthesis attribute INIT_0C of CH0_antialias_imdct_coefficient_RAM is "256'hC73BE272085A2B3C3E7B3B202263FD35D90AC2F63D09D90A02CA2263C4DF3E7B"
// Coe i = 6, k = 0-17
// synthesis attribute INIT_0D of CH0_antialias_imdct_coefficient_RAM is "256'h085A133ED4C33B20C00F38C4D90A0DDA133E32C63FF035FA187DF225D0D0C08C"
// Coe i = 24, k = 0-17
// synthesis attribute INIT_0E of CH0_antialias_imdct_coefficient_RAM is "256'h2F2F187DFD35E272CD39C184C18432C6E27202CA187DD0D03D09C08C35FADD9C"
// Coe i = 7, k = 0-17
// synthesis attribute INIT_0F of CH0_antialias_imdct_coefficient_RAM is "256'hCD3926F5E782085AF225D90AC73BC00FC4DFD4C3ECC1085A226335FA3F733D09"
// Coe i = 25, k = 0-17
// synthesis attribute INIT_10 of CH0_antialias_imdct_coefficient_RAM is "256'hC4DFC08C3F73C4DF32C6D90A187DF7A5F7A5187DD90A32C6C4DF3F73C08C3B20"
// synthesis attribute INIT_11 of CH0_antialias_imdct_coefficient_RAM is "256'h085A187D26F532C63B203F733F733B2032C626F5187D085AF7A5E782D90ACD39"
// Coe i = 8, k = 0-17
// synthesis attribute INIT_12 of CH0_antialias_imdct_coefficient_RAM is "256'hC1843D09C4DF38C4CA0532C6D0D02B3CD90A2263E272187DECC10DDAF7A502CA"
// Coe i = 26, k = 0-17
// synthesis attribute INIT_13 of CH0_antialias_imdct_coefficient_RAM is "256'hE782E272DD9CD90AD4C3D0D0CD39CA05C73BC4DFC2F6C184C08CC00FC00F3F73"
// Coe i = 9, k = 0-17
// synthesis attribute INIT_14 of CH0_antialias_imdct_coefficient_RAM is "256'h35FACD392F2FD4C326F5DD9C1D8DE782133EF225085AFD35FD35F7A5F225ECC1"
// Coe i = 27, k = 0-17
// synthesis attribute INIT_15 of CH0_antialias_imdct_coefficient_RAM is "256'hD4C3D0D0CD39CA05C73BC4DFC2F6C184C08CC00F3FF0C08C3E7BC2F63B20C73B"
// Coe i = 10, k = 0-17
// synthesis attribute INIT_16 of CH0_antialias_imdct_coefficient_RAM is "256'h3B20C08C3F73C4DF32C6D90A187DF7A5FD35F7A5F225ECC1E782E272DD9CD90A"
// Coe i = 28, k = 0-17
// synthesis attribute INIT_17 of CH0_antialias_imdct_coefficient_RAM is "256'hF7A5E782D90ACD39C4DFC08CC08C3B20CD3926F5E782085A085AE78226F5CD39"
// Coe i = 11, k = 0-17
// synthesis attribute INIT_18 of CH0_antialias_imdct_coefficient_RAM is "256'h3FF0C73B26F5F225085A187D26F532C63B203F733F733B2032C626F5187D085A"
// Coe i = 29, k = 0-17
// synthesis attribute INIT_19 of CH0_antialias_imdct_coefficient_RAM is "256'hCD39C1843E7BCD391D8DFD35E7822F2FC2F63F73CA052263F7A5ECC12B3CC4DF"
// synthesis attribute INIT_1A of CH0_antialias_imdct_coefficient_RAM is "256'hF225D90AC73BC00FC4DFD4C3ECC1085A226335FA3F733D092F2F187DFD35E272"
// Coe i = 12, k = 0-17
// synthesis attribute INIT_1B of CH0_antialias_imdct_coefficient_RAM is "256'hFD35DD9C3B20C1842B3CF7A5E27238C4C08C2F2FF225E78235FAC00F32C6ECC1"
// Coe i = 30, k = 0-17
// synthesis attribute INIT_1C of CH0_antialias_imdct_coefficient_RAM is "256'h187DF225D0D0C08CC73BE272085A2B3C3E7B3B202263FD35D90AC2F6C2F626F5"
// Coe i = 13, k = 0-17
// synthesis attribute INIT_1D of CH0_antialias_imdct_coefficient_RAM is "256'h187DC4DF3B20E782E7823B20C4DF187D187DC4DF3B20E782133E32C63FF035FA"
// Coe i = 31, k = 0-17
// synthesis attribute INIT_1E of CH0_antialias_imdct_coefficient_RAM is "256'hE782C4DFC4DFE782187D3B203B20187DE782C4DF3B20E782E7823B20C4DF187D"
// Coe i = 14, k = 0-17
// synthesis attribute INIT_1F of CH0_antialias_imdct_coefficient_RAM is "256'h32C602CACA053B20F225D4C33F73E272E782C4DFC4DFE782187D3B203B20187D"
// Coe i = 32, k = 0-17
// synthesis attribute INIT_20 of CH0_antialias_imdct_coefficient_RAM is "256'hDD9C187D3E7B2F2FF7A5C73BC73B085A2F2FC184187D2263C00F26F5133EC2F6"
// Coe i = 15, k = 0-17
// synthesis attribute INIT_21 of CH0_antialias_imdct_coefficient_RAM is "256'hD0D0ECC13F73DD9C1D8D3F732B3CF225C4DFCA05FD3532C63D09133ED90AC00F"
// Coe i = 33, k = 0-17
// synthesis attribute INIT_22 of CH0_antialias_imdct_coefficient_RAM is "256'h085ACA0535FA085AC2F62B3C187DC00F1D8D26F5C1840DDA32C6C73BFD353B20"
// synthesis attribute INIT_23 of CH0_antialias_imdct_coefficient_RAM is "256'hDD9CC08CECC12F2F3B2002CAC73BCD390DDA3E7B26F5E272C00FE7822B3C3D09"
// Coe i = 16, k = 0-17
// synthesis attribute INIT_24 of CH0_antialias_imdct_coefficient_RAM is "256'h3F73F7A5C4DF26F526F5C4DFF7A53F73E782CD3932C6187DC08C085A3B20D90A"
// Coe i = 34, k = 0-17
// synthesis attribute INIT_25 of CH0_antialias_imdct_coefficient_RAM is "256'hE78232C632C6E782C08CF7A53B2026F5D90AC4DF085A3F73187DCD39CD39E782"
// Coe i = 17, k = 0-17
// synthesis attribute INIT_26 of CH0_antialias_imdct_coefficient_RAM is "256'hC184F7A53FF0FD35C08C0DDA3D09E782C73B226332C6D4C326F53B20F7A5C08C"
// Coe i = 35, k = 0-17
// synthesis attribute INIT_27 of CH0_antialias_imdct_coefficient_RAM is "256'hFD35C00FF7A53E7B133EC4DFE27235FA26F5D0D02F2F26F5CA05E2723B20133E"
// Constant 0 (648-655)...
// synthesis attribute INIT_28 of CH0_antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000D4C3CD39226338C4E782C2F60DDA3F73"
// window coefficient for IMDCT block type 2 (656-667)...
// Constant 1 (668-703)...
// synthesis attribute INIT_29 of CH0_antialias_imdct_coefficient_RAM is "256'h4000400040004000085A187D26F532C63B203F733F733B2032C626F5187D085A"
// synthesis attribute INIT_2A of CH0_antialias_imdct_coefficient_RAM is "256'h4000400040004000400040004000400040004000400040004000400040004000"
// synthesis attribute INIT_2B of CH0_antialias_imdct_coefficient_RAM is "256'h4000400040004000400040004000400040004000400040004000400040004000"
// window coefficient for IMDCT block type 0 (704-767)...(index: 0, 18, 1, 19, 2, 20....)
// synthesis attribute INIT_2C of CH0_antialias_imdct_coefficient_RAM is "256'h32C626F535FA226338C41D8D3B20187D3D09133E3E7B0DDA3F73085A3FF002CA"
// synthesis attribute INIT_2D of CH0_antialias_imdct_coefficient_RAM is "256'h0DDA3E7B133E3D09187D3B201D8D38C4226335FA26F532C62B3C2F2F2F2F2B3C"
// Constant 0 (648-655)...
// synthesis attribute INIT_2E of CH0_antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000000000000000000002CA3FF0085A3F73"
// synthesis attribute INIT_2F of CH0_antialias_imdct_coefficient_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// window coefficient for IMDCT block type 1 (768-831)...(index: 0, 18, 1, 19, 2, 20....)
// synthesis attribute INIT_30 of CH0_antialias_imdct_coefficient_RAM is "256'h3B2026F53F73226340001D8D4000187D4000133E40000DDA4000085A400002CA"
// synthesis attribute INIT_31 of CH0_antialias_imdct_coefficient_RAM is "256'h00003E7B00003D0900003B20000038C4085A35FA187D32C626F52F2F32C62B3C"
// Constant 0 (648-655)...
// synthesis attribute INIT_32 of CH0_antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000000000000000000000003FF000003F73"
// synthesis attribute INIT_33 of CH0_antialias_imdct_coefficient_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// window coefficient for IMDCT block type 3 (832-895)...(index: 0, 18, 1, 19, 2, 20....)
// synthesis attribute INIT_34 of CH0_antialias_imdct_coefficient_RAM is "256'h32C6187D35FA085A38C400003B2000003D0900003E7B00003F7300003FF00000"
// synthesis attribute INIT_35 of CH0_antialias_imdct_coefficient_RAM is "256'h0DDA4000133E4000187D40001D8D400022633F7326F53B202B3C32C62F2F26F5"
// Constant 0 (648-655)...
// synthesis attribute INIT_36 of CH0_antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000000000000000000002CA4000085A4000"
// synthesis attribute INIT_37 of CH0_antialias_imdct_coefficient_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// COS coefficient for for IMDCT short block (896-967)...
// synthesis attribute INIT_38 of CH0_antialias_imdct_coefficient_RAM is "256'hCD3926F5E782085A3B20E782E7823B20C4DF187DCD39E7823F73F7A5C4DF26F5"
// synthesis attribute INIT_39 of CH0_antialias_imdct_coefficient_RAM is "256'h3B20D90AC4DF187D187DC4DF3B20E7823F73C4DF32C6D90A187DF7A5C08C3B20"
// synthesis attribute INIT_3A of CH0_antialias_imdct_coefficient_RAM is "256'h187D3B203B20187DE782C4DFD90AC4DF085A3F73187DCD3932C6187DC08C085A"
// synthesis attribute INIT_3B of CH0_antialias_imdct_coefficient_RAM is "256'h3B20187DE782C4DFF7A5E782D90ACD39C4DFC08CF7A5E782D90ACD39C4DFC08C"
// Constant -1 (968-999)...
// synthesis attribute INIT_3C of CH0_antialias_imdct_coefficient_RAM is "256'hC000C000C000C000C000C000C000C000D90AC4DF085A3F73187DCD39187D3B20"
// synthesis attribute INIT_3D of CH0_antialias_imdct_coefficient_RAM is "256'hC000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000"
// CS coefficient (1000-1007)...
// synthesis attribute INIT_3E of CH0_antialias_imdct_coefficient_RAM is "256'h3FFF3FFE3FF23FB63EEE3CC6386E36E1C000C000C000C000C000C000C000C000"
// CA coefficient (1008-1015)...
// -CA coefficient (1016-1023)...
// synthesis attribute INIT_3F of CH0_antialias_imdct_coefficient_RAM is "256'h003C00E8029F060D0BA4140E1E3020EDFFC3FF17FD60F9F2F45BEBF1E1CFDF12"

// synthesis translate_off

defparam CH0_antialias_imdct_coefficient_RAM.INIT_00 = 256'h35FA_1D8D_C4DF_ECC1_3E7B_085A_C00F_02CA_3F73_F225_C2F6_187D_38C4_DD9C_CD39_2B3C;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_01 = 256'hE782_C2F6_0DDA_3F73_FD35_C00F_F7A5_3E7B_133E_C4DF_E272_35FA_26F5_D0D0_D0D0_D90A;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_02 = 256'hD90A_3B20_085A_C08C_187D_32C6_CD39_E782_3F73_F7A5_C4DF_26F5_D4C3_CD39_2263_38C4;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_03 = 256'hC08C_F7A5_3B20_26F5_D90A_C4DF_085A_3F73_187D_CD39_32C6_187D_C08C_085A_3B20_D90A;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_04 = 256'hCD39_38C4_02CA_C4DF_2F2F_133E_C08C_2263_26F5_3B20_F7A5_C08C_E782_32C6_32C6_E782;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_05 = 256'hC00F_E782_2B3C_3D09_085A_CA05_CA05_F7A5_3D09_D4C3_E782_3FF0_E272_D90A_3E7B_F225;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_06 = 256'h0DDA_2B3C_C08C_1D8D_DD9C_C08C_ECC1_2F2F_3B20_02CA_C73B_CD39_0DDA_3E7B_26F5_E272;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_07 = 256'hF7A5_C73B_38C4_F7A5_D0D0_3E7B_E782_DD9C_3FF0_D90A_ECC1_3D09_CD39_FD35_35FA_C4DF;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_08 = 256'h1D8D_3F73_2B3C_F225_C4DF_CA05_FD35_32C6_3D09_133E_D90A_C00F_DD9C_187D_3E7B_2F2F;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_09 = 256'h187D_C4DF_3B20_E782_E782_3B20_C4DF_187D_187D_C4DF_3B20_E782_E782_3B20_C4DF_187D;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_0A = 256'h187D_3B20_3B20_187D_E782_C4DF_C4DF_E782_187D_3B20_3B20_187D_E782_C4DF_C4DF_187D;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_0B = 256'hD4C3_085A_1D8D_C73B_3F73_D0D0_0DDA_187D_CA05_3FF0_CD39_133E_E782_C4DF_C4DF_E782;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_0C = 256'hC73B_E272_085A_2B3C_3E7B_3B20_2263_FD35_D90A_C2F6_3D09_D90A_02CA_2263_C4DF_3E7B;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_0D = 256'h085A_133E_D4C3_3B20_C00F_38C4_D90A_0DDA_133E_32C6_3FF0_35FA_187D_F225_D0D0_C08C;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_0E = 256'h2F2F_187D_FD35_E272_CD39_C184_C184_32C6_E272_02CA_187D_D0D0_3D09_C08C_35FA_DD9C;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_0F = 256'hCD39_26F5_E782_085A_F225_D90A_C73B_C00F_C4DF_D4C3_ECC1_085A_2263_35FA_3F73_3D09;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_10 = 256'hC4DF_C08C_3F73_C4DF_32C6_D90A_187D_F7A5_F7A5_187D_D90A_32C6_C4DF_3F73_C08C_3B20;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_11 = 256'h085A_187D_26F5_32C6_3B20_3F73_3F73_3B20_32C6_26F5_187D_085A_F7A5_E782_D90A_CD39;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_12 = 256'hC184_3D09_C4DF_38C4_CA05_32C6_D0D0_2B3C_D90A_2263_E272_187D_ECC1_0DDA_F7A5_02CA;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_13 = 256'hE782_E272_DD9C_D90A_D4C3_D0D0_CD39_CA05_C73B_C4DF_C2F6_C184_C08C_C00F_C00F_3F73;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_14 = 256'h35FA_CD39_2F2F_D4C3_26F5_DD9C_1D8D_E782_133E_F225_085A_FD35_FD35_F7A5_F225_ECC1;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_15 = 256'hD4C3_D0D0_CD39_CA05_C73B_C4DF_C2F6_C184_C08C_C00F_3FF0_C08C_3E7B_C2F6_3B20_C73B;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_16 = 256'h3B20_C08C_3F73_C4DF_32C6_D90A_187D_F7A5_FD35_F7A5_F225_ECC1_E782_E272_DD9C_D90A;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_17 = 256'hF7A5_E782_D90A_CD39_C4DF_C08C_C08C_3B20_CD39_26F5_E782_085A_085A_E782_26F5_CD39;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_18 = 256'h3FF0_C73B_26F5_F225_085A_187D_26F5_32C6_3B20_3F73_3F73_3B20_32C6_26F5_187D_085A;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_19 = 256'hCD39_C184_3E7B_CD39_1D8D_FD35_E782_2F2F_C2F6_3F73_CA05_2263_F7A5_ECC1_2B3C_C4DF;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_1A = 256'hF225_D90A_C73B_C00F_C4DF_D4C3_ECC1_085A_2263_35FA_3F73_3D09_2F2F_187D_FD35_E272;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_1B = 256'hFD35_DD9C_3B20_C184_2B3C_F7A5_E272_38C4_C08C_2F2F_F225_E782_35FA_C00F_32C6_ECC1;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_1C = 256'h187D_F225_D0D0_C08C_C73B_E272_085A_2B3C_3E7B_3B20_2263_FD35_D90A_C2F6_C2F6_26F5;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_1D = 256'h187D_C4DF_3B20_E782_E782_3B20_C4DF_187D_187D_C4DF_3B20_E782_133E_32C6_3FF0_35FA;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_1E = 256'hE782_C4DF_C4DF_E782_187D_3B20_3B20_187D_E782_C4DF_3B20_E782_E782_3B20_C4DF_187D;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_1F = 256'h32C6_02CA_CA05_3B20_F225_D4C3_3F73_E272_E782_C4DF_C4DF_E782_187D_3B20_3B20_187D;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_20 = 256'hDD9C_187D_3E7B_2F2F_F7A5_C73B_C73B_085A_2F2F_C184_187D_2263_C00F_26F5_133E_C2F6;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_21 = 256'hD0D0_ECC1_3F73_DD9C_1D8D_3F73_2B3C_F225_C4DF_CA05_FD35_32C6_3D09_133E_D90A_C00F;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_22 = 256'h085A_CA05_35FA_085A_C2F6_2B3C_187D_C00F_1D8D_26F5_C184_0DDA_32C6_C73B_FD35_3B20;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_23 = 256'hDD9C_C08C_ECC1_2F2F_3B20_02CA_C73B_CD39_0DDA_3E7B_26F5_E272_C00F_E782_2B3C_3D09;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_24 = 256'h3F73_F7A5_C4DF_26F5_26F5_C4DF_F7A5_3F73_E782_CD39_32C6_187D_C08C_085A_3B20_D90A;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_25 = 256'hE782_32C6_32C6_E782_C08C_F7A5_3B20_26F5_D90A_C4DF_085A_3F73_187D_CD39_CD39_E782;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_26 = 256'hC184_F7A5_3FF0_FD35_C08C_0DDA_3D09_E782_C73B_2263_32C6_D4C3_26F5_3B20_F7A5_C08C;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_27 = 256'hFD35_C00F_F7A5_3E7B_133E_C4DF_E272_35FA_26F5_D0D0_2F2F_26F5_CA05_E272_3B20_133E;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_28 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_D4C3_CD39_2263_38C4_E782_C2F6_0DDA_3F73;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_29 = 256'h4000_4000_4000_4000_085A_187D_26F5_32C6_3B20_3F73_3F73_3B20_32C6_26F5_187D_085A;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_2A = 256'h4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_2B = 256'h4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_2C = 256'h32C6_26F5_35FA_2263_38C4_1D8D_3B20_187D_3D09_133E_3E7B_0DDA_3F73_085A_3FF0_02CA;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_2D = 256'h0DDA_3E7B_133E_3D09_187D_3B20_1D8D_38C4_2263_35FA_26F5_32C6_2B3C_2F2F_2F2F_2B3C;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_2E = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_02CA_3FF0_085A_3F73;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_2F = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_30 = 256'h3B20_26F5_3F73_2263_4000_1D8D_4000_187D_4000_133E_4000_0DDA_4000_085A_4000_02CA;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_31 = 256'h0000_3E7B_0000_3D09_0000_3B20_0000_38C4_085A_35FA_187D_32C6_26F5_2F2F_32C6_2B3C;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_32 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_3FF0_0000_3F73;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_33 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_34 = 256'h32C6_187D_35FA_085A_38C4_0000_3B20_0000_3D09_0000_3E7B_0000_3F73_0000_3FF0_0000;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_35 = 256'h0DDA_4000_133E_4000_187D_4000_1D8D_4000_2263_3F73_26F5_3B20_2B3C_32C6_2F2F_26F5;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_36 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_02CA_4000_085A_4000;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_37 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_38 = 256'hCD39_26F5_E782_085A_3B20_E782_E782_3B20_C4DF_187D_CD39_E782_3F73_F7A5_C4DF_26F5;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_39 = 256'h3B20_D90A_C4DF_187D_187D_C4DF_3B20_E782_3F73_C4DF_32C6_D90A_187D_F7A5_C08C_3B20;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_3A = 256'h187D_3B20_3B20_187D_E782_C4DF_D90A_C4DF_085A_3F73_187D_CD39_32C6_187D_C08C_085A;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_3B = 256'h3B20_187D_E782_C4DF_F7A5_E782_D90A_CD39_C4DF_C08C_F7A5_E782_D90A_CD39_C4DF_C08C;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_3C = 256'hC000_C000_C000_C000_C000_C000_C000_C000_D90A_C4DF_085A_3F73_187D_CD39_187D_3B20;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_3D = 256'hC000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_3E = 256'h3FFF_3FFE_3FF2_3FB6_3EEE_3CC6_386E_36E1_C000_C000_C000_C000_C000_C000_C000_C000;
defparam CH0_antialias_imdct_coefficient_RAM.INIT_3F = 256'h003C_00E8_029F_060D_0BA4_140E_1E30_20ED_FFC3_FF17_FD60_F9F2_F45B_EBF1_E1CF_DF12;

// synthesis translate_on

RAMB16_S18 CH1_antialias_imdct_coefficient_RAM (
	.DO(CH1_data_out),
	.DOP(),
	.ADDR(CH1_address),
	.CLK(clock),
	.DI(16'h0),
	.DIP(2'b00),
	.EN(CH1_mem_en),
	.SSR(1'b0),
	.WE(1'b0)
);

// COS coefficient for IMDCT for normal block (0-647)...
// Coe i = 0, k = 0-17
// synthesis attribute INIT_00 of CH1_antialias_imdct_coefficient_RAM is "256'h35FA1D8DC4DFECC13E7B085AC00F02CA3F73F225C2F6187D38C4DD9CCD392B3C"
// Coe i = 18, k = 0-17
// synthesis attribute INIT_01 of CH1_antialias_imdct_coefficient_RAM is "256'hE782C2F60DDA3F73FD35C00FF7A53E7B133EC4DFE27235FA26F5D0D0D0D0D90A"
// Coe i = 1, k = 0-17
// synthesis attribute INIT_02 of CH1_antialias_imdct_coefficient_RAM is "256'hD90A3B20085AC08C187D32C6CD39E7823F73F7A5C4DF26F5D4C3CD39226338C4"
// Coe i = 19, k = 0-17
// synthesis attribute INIT_03 of CH1_antialias_imdct_coefficient_RAM is "256'hC08CF7A53B2026F5D90AC4DF085A3F73187DCD3932C6187DC08C085A3B20D90A"
// Coe i = 2, k = 0-17
// synthesis attribute INIT_04 of CH1_antialias_imdct_coefficient_RAM is "256'hCD3938C402CAC4DF2F2F133EC08C226326F53B20F7A5C08CE78232C632C6E782"
// Coe i = 20, k = 0-17
// synthesis attribute INIT_05 of CH1_antialias_imdct_coefficient_RAM is "256'hC00FE7822B3C3D09085ACA05CA05F7A53D09D4C3E7823FF0E272D90A3E7BF225"
// Coe i = 3, k = 0-17
// synthesis attribute INIT_06 of CH1_antialias_imdct_coefficient_RAM is "256'h0DDA2B3CC08C1D8DDD9CC08CECC12F2F3B2002CAC73BCD390DDA3E7B26F5E272"
// Coe i = 21, k = 0-17
// synthesis attribute INIT_07 of CH1_antialias_imdct_coefficient_RAM is "256'hF7A5C73B38C4F7A5D0D03E7BE782DD9C3FF0D90AECC13D09CD39FD3535FAC4DF"
// synthesis attribute INIT_08 of CH1_antialias_imdct_coefficient_RAM is "256'h1D8D3F732B3CF225C4DFCA05FD3532C63D09133ED90AC00FDD9C187D3E7B2F2F"
// Coe i = 4, k = 0-17
// synthesis attribute INIT_09 of CH1_antialias_imdct_coefficient_RAM is "256'h187DC4DF3B20E782E7823B20C4DF187D187DC4DF3B20E782E7823B20C4DF187D"
// Coe i = 22, k = 0-17
// synthesis attribute INIT_0A of CH1_antialias_imdct_coefficient_RAM is "256'h187D3B203B20187DE782C4DFC4DFE782187D3B203B20187DE782C4DFC4DF187D"
// Coe i = 5, k = 0-17
// synthesis attribute INIT_0B of CH1_antialias_imdct_coefficient_RAM is "256'hD4C3085A1D8DC73B3F73D0D00DDA187DCA053FF0CD39133EE782C4DFC4DFE782"
// Coe i = 23, k = 0-17
// synthesis attribute INIT_0C of CH1_antialias_imdct_coefficient_RAM is "256'hC73BE272085A2B3C3E7B3B202263FD35D90AC2F63D09D90A02CA2263C4DF3E7B"
// Coe i = 6, k = 0-17
// synthesis attribute INIT_0D of CH1_antialias_imdct_coefficient_RAM is "256'h085A133ED4C33B20C00F38C4D90A0DDA133E32C63FF035FA187DF225D0D0C08C"
// Coe i = 24, k = 0-17
// synthesis attribute INIT_0E of CH1_antialias_imdct_coefficient_RAM is "256'h2F2F187DFD35E272CD39C184C18432C6E27202CA187DD0D03D09C08C35FADD9C"
// Coe i = 7, k = 0-17
// synthesis attribute INIT_0F of CH1_antialias_imdct_coefficient_RAM is "256'hCD3926F5E782085AF225D90AC73BC00FC4DFD4C3ECC1085A226335FA3F733D09"
// Coe i = 25, k = 0-17
// synthesis attribute INIT_10 of CH1_antialias_imdct_coefficient_RAM is "256'hC4DFC08C3F73C4DF32C6D90A187DF7A5F7A5187DD90A32C6C4DF3F73C08C3B20"
// synthesis attribute INIT_11 of CH1_antialias_imdct_coefficient_RAM is "256'h085A187D26F532C63B203F733F733B2032C626F5187D085AF7A5E782D90ACD39"
// Coe i = 8, k = 0-17
// synthesis attribute INIT_12 of CH1_antialias_imdct_coefficient_RAM is "256'hC1843D09C4DF38C4CA0532C6D0D02B3CD90A2263E272187DECC10DDAF7A502CA"
// Coe i = 26, k = 0-17
// synthesis attribute INIT_13 of CH1_antialias_imdct_coefficient_RAM is "256'hE782E272DD9CD90AD4C3D0D0CD39CA05C73BC4DFC2F6C184C08CC00FC00F3F73"
// Coe i = 9, k = 0-17
// synthesis attribute INIT_14 of CH1_antialias_imdct_coefficient_RAM is "256'h35FACD392F2FD4C326F5DD9C1D8DE782133EF225085AFD35FD35F7A5F225ECC1"
// Coe i = 27, k = 0-17
// synthesis attribute INIT_15 of CH1_antialias_imdct_coefficient_RAM is "256'hD4C3D0D0CD39CA05C73BC4DFC2F6C184C08CC00F3FF0C08C3E7BC2F63B20C73B"
// Coe i = 10, k = 0-17
// synthesis attribute INIT_16 of CH1_antialias_imdct_coefficient_RAM is "256'h3B20C08C3F73C4DF32C6D90A187DF7A5FD35F7A5F225ECC1E782E272DD9CD90A"
// Coe i = 28, k = 0-17
// synthesis attribute INIT_17 of CH1_antialias_imdct_coefficient_RAM is "256'hF7A5E782D90ACD39C4DFC08CC08C3B20CD3926F5E782085A085AE78226F5CD39"
// Coe i = 11, k = 0-17
// synthesis attribute INIT_18 of CH1_antialias_imdct_coefficient_RAM is "256'h3FF0C73B26F5F225085A187D26F532C63B203F733F733B2032C626F5187D085A"
// Coe i = 29, k = 0-17
// synthesis attribute INIT_19 of CH1_antialias_imdct_coefficient_RAM is "256'hCD39C1843E7BCD391D8DFD35E7822F2FC2F63F73CA052263F7A5ECC12B3CC4DF"
// synthesis attribute INIT_1A of CH1_antialias_imdct_coefficient_RAM is "256'hF225D90AC73BC00FC4DFD4C3ECC1085A226335FA3F733D092F2F187DFD35E272"
// Coe i = 12, k = 0-17
// synthesis attribute INIT_1B of CH1_antialias_imdct_coefficient_RAM is "256'hFD35DD9C3B20C1842B3CF7A5E27238C4C08C2F2FF225E78235FAC00F32C6ECC1"
// Coe i = 30, k = 0-17
// synthesis attribute INIT_1C of CH1_antialias_imdct_coefficient_RAM is "256'h187DF225D0D0C08CC73BE272085A2B3C3E7B3B202263FD35D90AC2F6C2F626F5"
// Coe i = 13, k = 0-17
// synthesis attribute INIT_1D of CH1_antialias_imdct_coefficient_RAM is "256'h187DC4DF3B20E782E7823B20C4DF187D187DC4DF3B20E782133E32C63FF035FA"
// Coe i = 31, k = 0-17
// synthesis attribute INIT_1E of CH1_antialias_imdct_coefficient_RAM is "256'hE782C4DFC4DFE782187D3B203B20187DE782C4DF3B20E782E7823B20C4DF187D"
// Coe i = 14, k = 0-17
// synthesis attribute INIT_1F of CH1_antialias_imdct_coefficient_RAM is "256'h32C602CACA053B20F225D4C33F73E272E782C4DFC4DFE782187D3B203B20187D"
// Coe i = 32, k = 0-17
// synthesis attribute INIT_20 of CH1_antialias_imdct_coefficient_RAM is "256'hDD9C187D3E7B2F2FF7A5C73BC73B085A2F2FC184187D2263C00F26F5133EC2F6"
// Coe i = 15, k = 0-17
// synthesis attribute INIT_21 of CH1_antialias_imdct_coefficient_RAM is "256'hD0D0ECC13F73DD9C1D8D3F732B3CF225C4DFCA05FD3532C63D09133ED90AC00F"
// Coe i = 33, k = 0-17
// synthesis attribute INIT_22 of CH1_antialias_imdct_coefficient_RAM is "256'h085ACA0535FA085AC2F62B3C187DC00F1D8D26F5C1840DDA32C6C73BFD353B20"
// synthesis attribute INIT_23 of CH1_antialias_imdct_coefficient_RAM is "256'hDD9CC08CECC12F2F3B2002CAC73BCD390DDA3E7B26F5E272C00FE7822B3C3D09"
// Coe i = 16, k = 0-17
// synthesis attribute INIT_24 of CH1_antialias_imdct_coefficient_RAM is "256'h3F73F7A5C4DF26F526F5C4DFF7A53F73E782CD3932C6187DC08C085A3B20D90A"
// Coe i = 34, k = 0-17
// synthesis attribute INIT_25 of CH1_antialias_imdct_coefficient_RAM is "256'hE78232C632C6E782C08CF7A53B2026F5D90AC4DF085A3F73187DCD39CD39E782"
// Coe i = 17, k = 0-17
// synthesis attribute INIT_26 of CH1_antialias_imdct_coefficient_RAM is "256'hC184F7A53FF0FD35C08C0DDA3D09E782C73B226332C6D4C326F53B20F7A5C08C"
// Coe i = 35, k = 0-17
// synthesis attribute INIT_27 of CH1_antialias_imdct_coefficient_RAM is "256'hFD35C00FF7A53E7B133EC4DFE27235FA26F5D0D02F2F26F5CA05E2723B20133E"
// Constant 0 (648-655)...
// synthesis attribute INIT_28 of CH1_antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000D4C3CD39226338C4E782C2F60DDA3F73"
// window coefficient for IMDCT block type 2 (656-667)...
// Constant 1 (668-703)...
// synthesis attribute INIT_29 of CH1_antialias_imdct_coefficient_RAM is "256'h4000400040004000085A187D26F532C63B203F733F733B2032C626F5187D085A"
// synthesis attribute INIT_2A of CH1_antialias_imdct_coefficient_RAM is "256'h4000400040004000400040004000400040004000400040004000400040004000"
// synthesis attribute INIT_2B of CH1_antialias_imdct_coefficient_RAM is "256'h4000400040004000400040004000400040004000400040004000400040004000"
// window coefficient for IMDCT block type 0 (704-767)...(index: 0, 18, 1, 19, 2, 20....)
// synthesis attribute INIT_2C of CH1_antialias_imdct_coefficient_RAM is "256'h32C626F535FA226338C41D8D3B20187D3D09133E3E7B0DDA3F73085A3FF002CA"
// synthesis attribute INIT_2D of CH1_antialias_imdct_coefficient_RAM is "256'h0DDA3E7B133E3D09187D3B201D8D38C4226335FA26F532C62B3C2F2F2F2F2B3C"
// Constant 0 (648-655)...
// synthesis attribute INIT_2E of CH1_antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000000000000000000002CA3FF0085A3F73"
// synthesis attribute INIT_2F of CH1_antialias_imdct_coefficient_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// window coefficient for IMDCT block type 1 (768-831)...(index: 0, 18, 1, 19, 2, 20....)
// synthesis attribute INIT_30 of CH1_antialias_imdct_coefficient_RAM is "256'h3B2026F53F73226340001D8D4000187D4000133E40000DDA4000085A400002CA"
// synthesis attribute INIT_31 of CH1_antialias_imdct_coefficient_RAM is "256'h00003E7B00003D0900003B20000038C4085A35FA187D32C626F52F2F32C62B3C"
// Constant 0 (648-655)...
// synthesis attribute INIT_32 of CH1_antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000000000000000000000003FF000003F73"
// synthesis attribute INIT_33 of CH1_antialias_imdct_coefficient_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// window coefficient for IMDCT block type 3 (832-895)...(index: 0, 18, 1, 19, 2, 20....)
// synthesis attribute INIT_34 of CH1_antialias_imdct_coefficient_RAM is "256'h32C6187D35FA085A38C400003B2000003D0900003E7B00003F7300003FF00000"
// synthesis attribute INIT_35 of CH1_antialias_imdct_coefficient_RAM is "256'h0DDA4000133E4000187D40001D8D400022633F7326F53B202B3C32C62F2F26F5"
// Constant 0 (648-655)...
// synthesis attribute INIT_36 of CH1_antialias_imdct_coefficient_RAM is "256'h00000000000000000000000000000000000000000000000002CA4000085A4000"
// synthesis attribute INIT_37 of CH1_antialias_imdct_coefficient_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// COS coefficient for for IMDCT short block (896-967)...
// synthesis attribute INIT_38 of CH1_antialias_imdct_coefficient_RAM is "256'hCD3926F5E782085A3B20E782E7823B20C4DF187DCD39E7823F73F7A5C4DF26F5"
// synthesis attribute INIT_39 of CH1_antialias_imdct_coefficient_RAM is "256'h3B20D90AC4DF187D187DC4DF3B20E7823F73C4DF32C6D90A187DF7A5C08C3B20"
// synthesis attribute INIT_3A of CH1_antialias_imdct_coefficient_RAM is "256'h187D3B203B20187DE782C4DFD90AC4DF085A3F73187DCD3932C6187DC08C085A"
// synthesis attribute INIT_3B of CH1_antialias_imdct_coefficient_RAM is "256'h3B20187DE782C4DFF7A5E782D90ACD39C4DFC08CF7A5E782D90ACD39C4DFC08C"
// Constant -1 (968-999)...
// synthesis attribute INIT_3C of CH1_antialias_imdct_coefficient_RAM is "256'hC000C000C000C000C000C000C000C000D90AC4DF085A3F73187DCD39187D3B20"
// synthesis attribute INIT_3D of CH1_antialias_imdct_coefficient_RAM is "256'hC000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000"
// CS coefficient (1000-1007)...
// synthesis attribute INIT_3E of CH1_antialias_imdct_coefficient_RAM is "256'h3FFF3FFE3FF23FB63EEE3CC6386E36E1C000C000C000C000C000C000C000C000"
// CA coefficient (1008-1015)...
// -CA coefficient (1016-1023)...
// synthesis attribute INIT_3F of CH1_antialias_imdct_coefficient_RAM is "256'h003C00E8029F060D0BA4140E1E3020EDFFC3FF17FD60F9F2F45BEBF1E1CFDF12"

// synthesis translate_off

defparam CH1_antialias_imdct_coefficient_RAM.INIT_00 = 256'h35FA_1D8D_C4DF_ECC1_3E7B_085A_C00F_02CA_3F73_F225_C2F6_187D_38C4_DD9C_CD39_2B3C;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_01 = 256'hE782_C2F6_0DDA_3F73_FD35_C00F_F7A5_3E7B_133E_C4DF_E272_35FA_26F5_D0D0_D0D0_D90A;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_02 = 256'hD90A_3B20_085A_C08C_187D_32C6_CD39_E782_3F73_F7A5_C4DF_26F5_D4C3_CD39_2263_38C4;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_03 = 256'hC08C_F7A5_3B20_26F5_D90A_C4DF_085A_3F73_187D_CD39_32C6_187D_C08C_085A_3B20_D90A;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_04 = 256'hCD39_38C4_02CA_C4DF_2F2F_133E_C08C_2263_26F5_3B20_F7A5_C08C_E782_32C6_32C6_E782;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_05 = 256'hC00F_E782_2B3C_3D09_085A_CA05_CA05_F7A5_3D09_D4C3_E782_3FF0_E272_D90A_3E7B_F225;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_06 = 256'h0DDA_2B3C_C08C_1D8D_DD9C_C08C_ECC1_2F2F_3B20_02CA_C73B_CD39_0DDA_3E7B_26F5_E272;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_07 = 256'hF7A5_C73B_38C4_F7A5_D0D0_3E7B_E782_DD9C_3FF0_D90A_ECC1_3D09_CD39_FD35_35FA_C4DF;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_08 = 256'h1D8D_3F73_2B3C_F225_C4DF_CA05_FD35_32C6_3D09_133E_D90A_C00F_DD9C_187D_3E7B_2F2F;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_09 = 256'h187D_C4DF_3B20_E782_E782_3B20_C4DF_187D_187D_C4DF_3B20_E782_E782_3B20_C4DF_187D;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_0A = 256'h187D_3B20_3B20_187D_E782_C4DF_C4DF_E782_187D_3B20_3B20_187D_E782_C4DF_C4DF_187D;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_0B = 256'hD4C3_085A_1D8D_C73B_3F73_D0D0_0DDA_187D_CA05_3FF0_CD39_133E_E782_C4DF_C4DF_E782;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_0C = 256'hC73B_E272_085A_2B3C_3E7B_3B20_2263_FD35_D90A_C2F6_3D09_D90A_02CA_2263_C4DF_3E7B;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_0D = 256'h085A_133E_D4C3_3B20_C00F_38C4_D90A_0DDA_133E_32C6_3FF0_35FA_187D_F225_D0D0_C08C;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_0E = 256'h2F2F_187D_FD35_E272_CD39_C184_C184_32C6_E272_02CA_187D_D0D0_3D09_C08C_35FA_DD9C;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_0F = 256'hCD39_26F5_E782_085A_F225_D90A_C73B_C00F_C4DF_D4C3_ECC1_085A_2263_35FA_3F73_3D09;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_10 = 256'hC4DF_C08C_3F73_C4DF_32C6_D90A_187D_F7A5_F7A5_187D_D90A_32C6_C4DF_3F73_C08C_3B20;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_11 = 256'h085A_187D_26F5_32C6_3B20_3F73_3F73_3B20_32C6_26F5_187D_085A_F7A5_E782_D90A_CD39;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_12 = 256'hC184_3D09_C4DF_38C4_CA05_32C6_D0D0_2B3C_D90A_2263_E272_187D_ECC1_0DDA_F7A5_02CA;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_13 = 256'hE782_E272_DD9C_D90A_D4C3_D0D0_CD39_CA05_C73B_C4DF_C2F6_C184_C08C_C00F_C00F_3F73;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_14 = 256'h35FA_CD39_2F2F_D4C3_26F5_DD9C_1D8D_E782_133E_F225_085A_FD35_FD35_F7A5_F225_ECC1;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_15 = 256'hD4C3_D0D0_CD39_CA05_C73B_C4DF_C2F6_C184_C08C_C00F_3FF0_C08C_3E7B_C2F6_3B20_C73B;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_16 = 256'h3B20_C08C_3F73_C4DF_32C6_D90A_187D_F7A5_FD35_F7A5_F225_ECC1_E782_E272_DD9C_D90A;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_17 = 256'hF7A5_E782_D90A_CD39_C4DF_C08C_C08C_3B20_CD39_26F5_E782_085A_085A_E782_26F5_CD39;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_18 = 256'h3FF0_C73B_26F5_F225_085A_187D_26F5_32C6_3B20_3F73_3F73_3B20_32C6_26F5_187D_085A;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_19 = 256'hCD39_C184_3E7B_CD39_1D8D_FD35_E782_2F2F_C2F6_3F73_CA05_2263_F7A5_ECC1_2B3C_C4DF;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_1A = 256'hF225_D90A_C73B_C00F_C4DF_D4C3_ECC1_085A_2263_35FA_3F73_3D09_2F2F_187D_FD35_E272;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_1B = 256'hFD35_DD9C_3B20_C184_2B3C_F7A5_E272_38C4_C08C_2F2F_F225_E782_35FA_C00F_32C6_ECC1;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_1C = 256'h187D_F225_D0D0_C08C_C73B_E272_085A_2B3C_3E7B_3B20_2263_FD35_D90A_C2F6_C2F6_26F5;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_1D = 256'h187D_C4DF_3B20_E782_E782_3B20_C4DF_187D_187D_C4DF_3B20_E782_133E_32C6_3FF0_35FA;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_1E = 256'hE782_C4DF_C4DF_E782_187D_3B20_3B20_187D_E782_C4DF_3B20_E782_E782_3B20_C4DF_187D;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_1F = 256'h32C6_02CA_CA05_3B20_F225_D4C3_3F73_E272_E782_C4DF_C4DF_E782_187D_3B20_3B20_187D;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_20 = 256'hDD9C_187D_3E7B_2F2F_F7A5_C73B_C73B_085A_2F2F_C184_187D_2263_C00F_26F5_133E_C2F6;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_21 = 256'hD0D0_ECC1_3F73_DD9C_1D8D_3F73_2B3C_F225_C4DF_CA05_FD35_32C6_3D09_133E_D90A_C00F;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_22 = 256'h085A_CA05_35FA_085A_C2F6_2B3C_187D_C00F_1D8D_26F5_C184_0DDA_32C6_C73B_FD35_3B20;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_23 = 256'hDD9C_C08C_ECC1_2F2F_3B20_02CA_C73B_CD39_0DDA_3E7B_26F5_E272_C00F_E782_2B3C_3D09;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_24 = 256'h3F73_F7A5_C4DF_26F5_26F5_C4DF_F7A5_3F73_E782_CD39_32C6_187D_C08C_085A_3B20_D90A;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_25 = 256'hE782_32C6_32C6_E782_C08C_F7A5_3B20_26F5_D90A_C4DF_085A_3F73_187D_CD39_CD39_E782;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_26 = 256'hC184_F7A5_3FF0_FD35_C08C_0DDA_3D09_E782_C73B_2263_32C6_D4C3_26F5_3B20_F7A5_C08C;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_27 = 256'hFD35_C00F_F7A5_3E7B_133E_C4DF_E272_35FA_26F5_D0D0_2F2F_26F5_CA05_E272_3B20_133E;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_28 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_D4C3_CD39_2263_38C4_E782_C2F6_0DDA_3F73;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_29 = 256'h4000_4000_4000_4000_085A_187D_26F5_32C6_3B20_3F73_3F73_3B20_32C6_26F5_187D_085A;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_2A = 256'h4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_2B = 256'h4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000_4000;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_2C = 256'h32C6_26F5_35FA_2263_38C4_1D8D_3B20_187D_3D09_133E_3E7B_0DDA_3F73_085A_3FF0_02CA;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_2D = 256'h0DDA_3E7B_133E_3D09_187D_3B20_1D8D_38C4_2263_35FA_26F5_32C6_2B3C_2F2F_2F2F_2B3C;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_2E = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_02CA_3FF0_085A_3F73;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_2F = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_30 = 256'h3B20_26F5_3F73_2263_4000_1D8D_4000_187D_4000_133E_4000_0DDA_4000_085A_4000_02CA;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_31 = 256'h0000_3E7B_0000_3D09_0000_3B20_0000_38C4_085A_35FA_187D_32C6_26F5_2F2F_32C6_2B3C;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_32 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_3FF0_0000_3F73;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_33 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_34 = 256'h32C6_187D_35FA_085A_38C4_0000_3B20_0000_3D09_0000_3E7B_0000_3F73_0000_3FF0_0000;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_35 = 256'h0DDA_4000_133E_4000_187D_4000_1D8D_4000_2263_3F73_26F5_3B20_2B3C_32C6_2F2F_26F5;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_36 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_02CA_4000_085A_4000;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_37 = 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_38 = 256'hCD39_26F5_E782_085A_3B20_E782_E782_3B20_C4DF_187D_CD39_E782_3F73_F7A5_C4DF_26F5;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_39 = 256'h3B20_D90A_C4DF_187D_187D_C4DF_3B20_E782_3F73_C4DF_32C6_D90A_187D_F7A5_C08C_3B20;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_3A = 256'h187D_3B20_3B20_187D_E782_C4DF_D90A_C4DF_085A_3F73_187D_CD39_32C6_187D_C08C_085A;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_3B = 256'h3B20_187D_E782_C4DF_F7A5_E782_D90A_CD39_C4DF_C08C_F7A5_E782_D90A_CD39_C4DF_C08C;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_3C = 256'hC000_C000_C000_C000_C000_C000_C000_C000_D90A_C4DF_085A_3F73_187D_CD39_187D_3B20;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_3D = 256'hC000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000_C000;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_3E = 256'h3FFF_3FFE_3FF2_3FB6_3EEE_3CC6_386E_36E1_C000_C000_C000_C000_C000_C000_C000_C000;
defparam CH1_antialias_imdct_coefficient_RAM.INIT_3F = 256'h003C_00E8_029F_060D_0BA4_140E_1E30_20ED_FFC3_FF17_FD60_F9F2_F45B_EBF1_E1CF_DF12;

// synthesis translate_on
*/
endmodule
