// 
//  MAC_MP3: A Low Energy Implementation of an Audio Decoder
//
//  Copyright (C) 2007 McMaster University
// 
//==============================================================================
// 
// This file is part of MAC_MP3
// 
// MAC_MP3 is distributed in the hope that it will be useful for further research,
// but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY
// or FITNESS FOR A PARTICULAR PURPOSE. MAC_MP3 is free; you can redistribute it
// and/or modify it provided that proper reference is provided to the authors. See
// the documents included in the "doc" folder for further details.
//
//==============================================================================


`timescale 1ns / 100ps

module bigrom(clk,addressA,dataoutA,addressB,dataoutB);
  input clk;
  input [14:0] addressA;
  output [15:0] dataoutA;
  input [14:0] addressB;
  output [15:0] dataoutB;

  reg [4:0] addrmuxA;
  reg [4:0] addrmuxB;
  //wire addrmuxA;
  //wire addrmuxB;
  wire [15:0] memdataA [31:0];
  wire [15:0] memdataB [31:0];
  
  //assign addrmuxA = addressA[10];
  //assign addrmuxB = addressB[10];
  assign dataoutA = memdataA[addrmuxA];
  assign dataoutB = memdataB[addrmuxB];
  
  always @ (posedge clk)
  begin
    addrmuxA <= addressA[14:10];
    addrmuxB <= addressB[14:10];
  end
  
  RAMB16_S18_S18 bigblock0 (
    .DOA(memdataA[0]),
    .DOB(memdataB[0]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );
  
  RAMB16_S18_S18 bigblock1 (
    .DOA(memdataA[1]),
    .DOB(memdataB[1]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock2 (
    .DOA(memdataA[2]),
    .DOB(memdataB[2]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock3 (
    .DOA(memdataA[3]),
    .DOB(memdataB[3]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock4 (
    .DOA(memdataA[4]),
    .DOB(memdataB[4]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock5 (
    .DOA(memdataA[5]),
    .DOB(memdataB[5]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock6 (
    .DOA(memdataA[6]),
    .DOB(memdataB[6]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock7 (
    .DOA(memdataA[7]),
    .DOB(memdataB[7]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock8 (
    .DOA(memdataA[8]),
    .DOB(memdataB[8]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock9 (
    .DOA(memdataA[9]),
    .DOB(memdataB[9]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblockA (
    .DOA(memdataA[5'hA]),
    .DOB(memdataB[5'hA]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblockB (
    .DOA(memdataA[5'hB]),
    .DOB(memdataB[5'hB]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblockC (
    .DOA(memdataA[5'hC]),
    .DOB(memdataB[5'hC]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblockD (
    .DOA(memdataA[5'hD]),
    .DOB(memdataB[5'hD]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblockE (
    .DOA(memdataA[5'hE]),
    .DOB(memdataB[5'hE]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblockF (
    .DOA(memdataA[5'hF]),
    .DOB(memdataB[5'hF]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock10 (
    .DOA(memdataA[5'h10]),
    .DOB(memdataB[5'h10]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock11 (
    .DOA(memdataA[5'h11]),
    .DOB(memdataB[5'h11]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock12 (
    .DOA(memdataA[5'h12]),
    .DOB(memdataB[5'h12]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock13 (
    .DOA(memdataA[5'h13]),
    .DOB(memdataB[5'h13]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock14 (
    .DOA(memdataA[5'h14]),
    .DOB(memdataB[5'h14]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock15 (
    .DOA(memdataA[5'h15]),
    .DOB(memdataB[5'h15]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock16 (
    .DOA(memdataA[5'h16]),
    .DOB(memdataB[5'h16]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock17 (
    .DOA(memdataA[5'h17]),
    .DOB(memdataB[5'h17]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock18 (
    .DOA(memdataA[5'h18]),
    .DOB(memdataB[5'h18]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock19 (
    .DOA(memdataA[5'h19]),
    .DOB(memdataB[5'h19]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock1A (
    .DOA(memdataA[5'h1A]),
    .DOB(memdataB[5'h1A]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock1B (
    .DOA(memdataA[5'h1B]),
    .DOB(memdataB[5'h1B]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock1C(
    .DOA(memdataA[5'h1C]),
    .DOB(memdataB[5'h1C]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock1D (
    .DOA(memdataA[5'h1D]),
    .DOB(memdataB[5'h1D]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock1E (
    .DOA(memdataA[5'h1E]),
    .DOB(memdataB[5'h1E]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  RAMB16_S18_S18 bigblock1F (
    .DOA(memdataA[5'h1F]),
    .DOB(memdataB[5'h1F]),
    .DOPA(),
    .DOPB(),
    .ADDRA(addressA[9:0]),
    .ADDRB(addressB[9:0]),
    .CLKA(clk),
    .CLKB(clk),
    .DIA(16'h0000),
    .DIB(16'h0000),
    .DIPA(2'b00),
    .DIPB(2'b00),
    .ENA(1'b1),
    .ENB(1'b1),
    .SSRA(1'b0),
    .SSRB(1'b0),
    .WEA(1'b0),
    .WEB(1'b0)
  );

  `include "./rom/mp3_src.v"
//  `include "memory/rom/06.v"
  //`include "memory/rom/nissin.v"
  //`include "memory/rom/Pancakes.v"
  //`include "memory/rom/McDonaldSummer.v"
  //`include "memory/rom/funky.v"
  ////`include "memory/rom/part_of_me.v"
  //`include "memory/rom/spot2.v"
  //`include "memory/rom/spot3.v"
  //`include "memory/rom/plane.v"
  //`include "memory/rom/KillBill.v"
  //`include "memory/rom/beer.v"
  //`include "memory/rom/beer1.v"

// spot1.v
/*  
// synthesis attribute INIT_00 of bigblock0 is "256'h82ed003df1806b1c08610005c61c2b5f30a30400ee3e4eda04d604807274fffb"
// synthesis attribute INIT_01 of bigblock0 is "256'h7343a791b2859e3ca4a0811d1c98358b8a48bb10a602e15255c6061b00006b86"
// synthesis attribute INIT_02 of bigblock0 is "256'hf566d4be836d202b7f0868e1aaa89aa80cbebe541a80d1c3b949b60c8bc22354"
// synthesis attribute INIT_03 of bigblock0 is "256'hb84e1b5cf51ae993f3b60d185f24e93eb87ca8d0541234b3ab51a44a543ce398"
// synthesis attribute INIT_04 of bigblock0 is "256'ha2aace9a2a1be26f1d32e40d9a052b3abb9b89e5892426260ac664ccd523267c"
// synthesis attribute INIT_05 of bigblock0 is "256'h9ffe01dc140201c0c01ce57c34f151dc84267d447186f406ca444d66bacc28a0"
// synthesis attribute INIT_06 of bigblock0 is "256'he79e148a21bf04401d257933edc12b4fea720674d632db4783036db2b6dbdb6d"
// synthesis attribute INIT_07 of bigblock0 is "256'hc5d713590184c7bfef7c1aa3cc78df40baf1e3050af10400e0001b07c68896f3"
// synthesis attribute INIT_08 of bigblock0 is "256'h905bbd0b114c84e65f786d83492400ee40000fe91b4160c62385b3e1cc88e8e1"
// synthesis attribute INIT_09 of bigblock0 is "256'h0e007274fffb3722907f6cc6445ca899bf8722cc40e4a32b012770ab4a2e9020"
// synthesis attribute INIT_0A of bigblock0 is "256'h7ad18c11245184ae2848a0db71a4755b304f0c42cb8a126040785126265c02d7"
// synthesis attribute INIT_0B of bigblock0 is "256'h705dbbd521040940a090e631d5ece5d45154753152a13bc5b5cf420882972699"
// synthesis attribute INIT_0C of bigblock0 is "256'hb05cfe22fd48c4197d88392639acb1747904b410a308d1e06cd8b84e516d8932"
// synthesis attribute INIT_0D of bigblock0 is "256'h8a9b680872238b809b8300000a20002336c2fc71d4ad8410c3abc4f424889249"
// synthesis attribute INIT_0E of bigblock0 is "256'h6cefbe2d95dca5e43892acbdf1ac4cc19131c3679e24411bb520d054031884b9"
// synthesis attribute INIT_0F of bigblock0 is "256'h162e8b0ad12faeb96aaa9289b48e44679b6a974ad2afb65844bcd8fa4abd58cb"
// synthesis attribute INIT_10 of bigblock0 is "256'h487b0802cbc12922e3cf1689284362d3047263389b907e824398345c58a55848"
// synthesis attribute INIT_11 of bigblock0 is "256'hd9233341fe6a0b51159164cc4350852cffff463fc840dad9e19c2468914bc2a6"
// synthesis attribute INIT_12 of bigblock0 is "256'h6b68fae5b36e28e476c2037ba45922832115a20a03074078330c4e47502951a6"
// synthesis attribute INIT_13 of bigblock0 is "256'he92359de03381b807274fffb6fe9ddcdaa5d94b39988da759665dc291939462c"
// synthesis attribute INIT_14 of bigblock0 is "256'h4c86337b846bc9088c81741407efe07198697ba44947120c0502bbdc17812dc8"
// synthesis attribute INIT_15 of bigblock0 is "256'h6665cace8eedea3163191e46fee4a18ecf621a543151373ba1462d74c2d11851"
// synthesis attribute INIT_16 of bigblock0 is "256'h08d48a39c1018f26409aeecd17403304fb05bfffdb4921d2663b69abc99cb95d"
// synthesis attribute INIT_17 of bigblock0 is "256'he418922d95e48918bb6f48fe6d02d178708107e437a110b70ba8448294d40c44"
// synthesis attribute INIT_18 of bigblock0 is "256'h41c24629de98ce6705faca792891bbcab320456b3952d126a1fa0516114d04ad"
// synthesis attribute INIT_19 of bigblock0 is "256'hf0850b2a71545841462ae67af485690bee5e6dd75e12b5943274f87f3cf75c05"
// synthesis attribute INIT_1A of bigblock0 is "256'h2410890ca1438f0f07809a338f2f7822344859dccf30b6d9e36d6536010049a4"
// synthesis attribute INIT_1B of bigblock0 is "256'h5c223b4d4fbc3ccb892c962d9761c0eb98d2e2945683a8acdba83b683a004b6a"
// synthesis attribute INIT_1C of bigblock0 is "256'h3ea37bff379dad7d489154af964f1b91c63a36fcfdf8cd2531f2d39b168ff1c8"
// synthesis attribute INIT_1D of bigblock0 is "256'h9bca18021e48612648de032528007074fffbed47f1a76c296f961dfed422357a"
// synthesis attribute INIT_1E of bigblock0 is "256'hf174e233cabd6431dff6b7d60c9d8468241104efe059187178c3651b344b0462"
// synthesis attribute INIT_1F of bigblock0 is "256'hc21187e6ee9515f9ab9182a55ca198ab781a6d86b91bb2a9fc00b52b5d513114"
// synthesis attribute INIT_20 of bigblock0 is "256'he7efb2ab5acaf870ca6563460de818df8b4b74aed864736ec414f9d23c48a100"
// synthesis attribute INIT_21 of bigblock0 is "256'h854c14686ea1956e3be58a2db0a65e1b12e5927128b9bd101a9dbb33f9add8c1"
// synthesis attribute INIT_22 of bigblock0 is "256'hff261bff400890a405089fe41e55c18b8806174e2c11cbcbb87d653253d7e320"
// synthesis attribute INIT_23 of bigblock0 is "256'h056f84df32213f440916008b2d809901ca994f892c8b86872575732ade9b9f01"
// synthesis attribute INIT_24 of bigblock0 is "256'hb79d63def3842c7d87cc71f2f8cf66ceef633b6895658e3964d0dc9033cf234d"
// synthesis attribute INIT_25 of bigblock0 is "256'hc4a45ce785c569b2768f9b82c2874143ac44309496b276e09db92738d079f197"
// synthesis attribute INIT_26 of bigblock0 is "256'h40130100d680d3a9c19c23db60d2b162a38112937fe6afa9f78d2fb28d92cec4"
// synthesis attribute INIT_27 of bigblock0 is "256'hfd774b040302bc04a13b881623375dc95c488003743bfb72f3ffe92c92567fff"
// synthesis attribute INIT_28 of bigblock0 is "256'h2489e82f000254c9e801be00d33a6d5eb7d524bf0808200c2ee44f0567c04498"
// synthesis attribute INIT_29 of bigblock0 is "256'h74e7c10e8935c1f18149eb2c5b24b2b4b8d94e35d21001f08c83e0b667971a4a"
// synthesis attribute INIT_2A of bigblock0 is "256'h1e26a6bc508d15ceff21e949d8f3ff3ca23bdd56a4dfec21752cd0489a9e9d48"
// synthesis attribute INIT_2B of bigblock0 is "256'h133db1edc6edeb9ca446ee8cfff041afe0116b622f3e73cdca637f8303d02506"
// synthesis attribute INIT_2C of bigblock0 is "256'h6a1b3aefa9eec57948baad41412213a285642a1012a700293640094926ba6a94"
// synthesis attribute INIT_2D of bigblock0 is "256'hd7bb90020f95fff7289e7ceb437dcbec3ccc518e8655912ac6c44e2b674ee8a9"
// synthesis attribute INIT_2E of bigblock0 is "256'h9bba472274ab0b34ca0313d01505b4bb2dab8cf5219ebba0885d14a8d699cc14"
// synthesis attribute INIT_2F of bigblock0 is "256'h04d3c151b8c67dfbb677b5a1cb7144ac3896b1a0d69abffe10414a406ea85073"
// synthesis attribute INIT_30 of bigblock0 is "256'h0c529c45297bd08ad265c8fc2709a5f8b0adacf510d7844d89a3b4d3012a0990"
// synthesis attribute INIT_31 of bigblock0 is "256'h67046f40a62427754c612340ac20a13bb0188615dd690d3f8003744ffb7204ff"
// synthesis attribute INIT_32 of bigblock0 is "256'hd6ab523fa91fe1458f0a9e604770ffbfe4c42efeab66841181bc803d348ceeb0"
// synthesis attribute INIT_33 of bigblock0 is "256'h0db1f5ec8e6511dbd965df4ce5eecd6154a4174fdab71d4da4fa6998ebd3655c"
// synthesis attribute INIT_34 of bigblock0 is "256'hb25d6801660854d18c1f54a4e58ba7610a01d41108cafffe892b5510a6401ba2"
// synthesis attribute INIT_35 of bigblock0 is "256'ha926045523efba904f18c3e6af0a222daa35bc8c2aaea2a1a9652ead00fc0cc8"
// synthesis attribute INIT_36 of bigblock0 is "256'h5feee7fa5e4e2a8e11c862a338bc0b29f4af27df9efb43fdfc67c4ebfc98295b"
// synthesis attribute INIT_37 of bigblock0 is "256'h2be097f6d4718696c01909301532973820f6718bc82ce2a15652a1b181f2db30"
// synthesis attribute INIT_38 of bigblock0 is "256'h1520080088b33a017ca470e846d128bb7e5d7e87c3391c290e48b0c26fffa046"
// synthesis attribute INIT_39 of bigblock0 is "256'h85d25ea30f6d8b7f1637f797303b12936c2cb890e28962e997700e2a9dcd4399"
// synthesis attribute INIT_3A of bigblock0 is "256'h745ffb724cff06ce3b424d2e00e4cf0661558412a8e121d1534ff3bac0b4242c"
// synthesis attribute INIT_3B of bigblock0 is "256'h810c248c6ea46d0a6bc0a7a403754c6d2374a90c229ba01887335d6112340003"
// synthesis attribute INIT_3C of bigblock0 is "256'h491e90ce925a8600b7ae6e48aa8a4674c0ddececfb76a7fe934ef334e558da48"
// synthesis attribute INIT_3D of bigblock0 is "256'hd24042526554a3ea02c251aabe9585317cf5dc0caa6215cc9c660f56fffb1d4a"
// synthesis attribute INIT_3E of bigblock0 is "256'hd38da0a85736af35ad8990c851f0d1bdacb6ea637b15b42e8dc833551f2c014b"
// synthesis attribute INIT_3F of bigblock0 is "256'hab322b6ff3dd673bd7d092a22c7d2b5190bada40d56bd5552235846682acec2e"
// synthesis attribute INIT_00 of bigblock1 is "256'hd634e6c7fffd24b7851860596b569dec774a40f88300ef4347b1c2c156540d7b"
// synthesis attribute INIT_01 of bigblock1 is "256'h2c91b674a9c82995001ab1f010128a4038ad20b1213b0625931f163c5369b1d3"
// synthesis attribute INIT_02 of bigblock1 is "256'hcc7a42bec111bce5819863ca6c2887a865cdd8ca134f6c63c88ce4415cb0be1b"
// synthesis attribute INIT_03 of bigblock1 is "256'h8b46377e05c3667171d0d191c1aa09b03eae9909d631c458b324813040626184"
// synthesis attribute INIT_04 of bigblock1 is "256'h5e69de3d8002746dfb7000ffa0396be176f168d57533cc38a30e2b9f3599a544"
// synthesis attribute INIT_05 of bigblock1 is "256'h6db226db1272980013156f34758a6d2083241f794c552234cc18429bf01be929"
// synthesis attribute INIT_06 of bigblock1 is "256'hb02918578000713a8464cb284619c07349483dfade067e0b94bf078647a919e4"
// synthesis attribute INIT_07 of bigblock1 is "256'hfbfbf71b90ead3596f45c73e46d15354df0facf50871307aac363094d56aa2ec"
// synthesis attribute INIT_08 of bigblock1 is "256'hb2acb7470523eee2dce88569e32ea33534a24e3dc5a528e1a63851ece7cc14de"
// synthesis attribute INIT_09 of bigblock1 is "256'hd9886db6c76b022cfda09ad7a6b510265f2c60aa3053a170203af9272d63b7ba"
// synthesis attribute INIT_0A of bigblock1 is "256'h50a641bb51390001e471282c96924e33427b8d2b85165cdb3958e0c27a5287ba"
// synthesis attribute INIT_0B of bigblock1 is "256'hec5bc25bd76b24a323d81ef0be4ca4d191fde706acab903f0483488675639dd7"
// synthesis attribute INIT_0C of bigblock1 is "256'h3e8aa8c62dad0efce5b6b265778fba515cd4dc11983339f160b70ab447d79cf6"
// synthesis attribute INIT_0D of bigblock1 is "256'h25e5a2b5c3cddb6c55b638ed40682cd01eb3886138d85010f87c0ea488964583"
// synthesis attribute INIT_0E of bigblock1 is "256'hdbed1c222b6868c9445f030e7c807274fffb409e1cc50472284c4388c13d0b21"
// synthesis attribute INIT_0F of bigblock1 is "256'hf654cf8138b2880551b4121345320d49b41389ef6074a46f7da5e10f740b0826"
// synthesis attribute INIT_10 of bigblock1 is "256'hc0d19dfd6306c730f3a3fb5392c9ab4cd8a4d627c36031605ae58af098a21718"
// synthesis attribute INIT_11 of bigblock1 is "256'h68d76d697b5dd6e8b96eb6034a9e1fe8c76ac49656d116e5b50f6ed477ddcbcb"
// synthesis attribute INIT_12 of bigblock1 is "256'ha106dc22a6e62e8efab257ff094e2a04b4ff5aeb7eae0397820d5705a8517335"
// synthesis attribute INIT_13 of bigblock1 is "256'h91691f79d2cdeeb931f13469222d033eaf00ae3dbf13c5c1b2160110c813be82"
// synthesis attribute INIT_14 of bigblock1 is "256'h9214fdedf682fe8bfc881f75834558c20e19a745ce21fa15f5a77ec0284ca4b3"
// synthesis attribute INIT_15 of bigblock1 is "256'h255936fc7e6bcab1b37e8f7da23f6f0ff3f09e5e25216a9d75ba0c5944f8c76d"
// synthesis attribute INIT_16 of bigblock1 is "256'h8f8006b54de169a4b441fe5197ff82828124a14421dd2d94815a65b8ebf8bde1"
// synthesis attribute INIT_17 of bigblock1 is "256'he0c824fc1f9c04cd61f397001c89a865000004048ad0846535e9f19f2bc69049"
// synthesis attribute INIT_18 of bigblock1 is "256'h511d704c0c43fbbc1bc11450e986485d02e88a807274fffb2fe77864e0e6b69a"
// synthesis attribute INIT_19 of bigblock1 is "256'h5fb8ebb189ccfa673dfcca67a27d1c031f24f58e0d88f0110b6ea06b20d67726"
// synthesis attribute INIT_1A of bigblock1 is "256'hde500786148436cb9355da9da7b1820e6e5c9af9fb9d3ba95d667ceb3606363a"
// synthesis attribute INIT_1B of bigblock1 is "256'he55e9065d96315400437d4a3b1625fff390133f7e755bbde1322d1020b35030b"
// synthesis attribute INIT_1C of bigblock1 is "256'hf363e0ca60cbc68e32afc1a625857a240297600083115a40c30077c6909a285e"
// synthesis attribute INIT_1D of bigblock1 is "256'h7c4eed36923b957637fb6e5c6cf7563103e5a66524864d3a2fb9e292f152928a"
// synthesis attribute INIT_1E of bigblock1 is "256'hca315e6d4404596cf044b90f335c9c5b7ac6bb71c36f8840ee3910e67dfc1582"
// synthesis attribute INIT_1F of bigblock1 is "256'h8eca8dcc0996e0ab305868613695fff8221700b3b6313c584b182753f9cc787e"
// synthesis attribute INIT_20 of bigblock1 is "256'h20cce2f524e02023fc78842c9a8d0220469ad1518000997684897647b50933fa"
// synthesis attribute INIT_21 of bigblock1 is "256'h61de52d865b498abb432ef719b52d6d7bc5572a285d1529e7836221b2029eac3"
// synthesis attribute INIT_22 of bigblock1 is "256'hc06a246d71a69cf9604c0c25db891a4114606926415c03029a807274fffb61f0"
// synthesis attribute INIT_23 of bigblock1 is "256'h42d8beb8b3ba99e8d5a18faa9da4d07dcb928da3fa5a5cc9f35c883024218b6e"
// synthesis attribute INIT_24 of bigblock1 is "256'h5a745839e496c640f68f95ff22e427fc21d4cd8b4282b69d52e709be4a1d3450"
// synthesis attribute INIT_25 of bigblock1 is "256'h8822848253729d3e4ebbbca9026f741e0013a24d00222d0975cb1a2a4596f49f"
// synthesis attribute INIT_26 of bigblock1 is "256'h718ff7e9d0a0651fa53dd8a6a7ff27127cc22291c438c1a4ebb1900fda8fe263"
// synthesis attribute INIT_27 of bigblock1 is "256'hb9439be6f02972a37f4e41272aa253042659f48d84a549923f2d4fcfc96731fc"
// synthesis attribute INIT_28 of bigblock1 is "256'hb3a82e458f767e81e7da428289da52b3f65545ff8828e8ac575fe292faefdcad"
// synthesis attribute INIT_29 of bigblock1 is "256'h542289ab71093fc119e43a7be624109384678b395c23d3c6cf33000019104728"
// synthesis attribute INIT_2A of bigblock1 is "256'h69dc9d5504139ea93cba6b884969b8cb4953aa199efcc9301024536afb1716e5"
// synthesis attribute INIT_2B of bigblock1 is "256'h7074fffbee4551b585416135a5ed82e42ed4e2abc903ceb86c05c0ec45db6d7d"
// synthesis attribute INIT_2C of bigblock1 is "256'h88c9a460872ec859987275a41925500c0c43dba91741430848c7445d0335a880"
// synthesis attribute INIT_2D of bigblock1 is "256'ha6ad70c4eb73632907c88957000fee8bbb92e34d00060600f68fc6ac12602fa8"
// synthesis attribute INIT_2E of bigblock1 is "256'h7367d23c5bf77328355c3301d86ba88d2953240dcfdc655d000b000554395244"
// synthesis attribute INIT_2F of bigblock1 is "256'h8bf0d7c2e396885b7673bbba2c29cbfe1f0a5be0699d126a8fb0a24b72156069"
// synthesis attribute INIT_30 of bigblock1 is "256'h5438ba7b2ab44abafc075e4f3ffab9d4eafa3f3343bf270f8b29e29d07c6b6d2"
// synthesis attribute INIT_31 of bigblock1 is "256'h480500c0cbea2b8ed7309f45a2338272fe9a72a8682e17cefbf5015f10a0ad3a"
// synthesis attribute INIT_32 of bigblock1 is "256'hda00d8194a566b9e16b2938c3cf5377e48683aeeca9ae17650f767b33f1a7880"
// synthesis attribute INIT_33 of bigblock1 is "256'h1f5346dfa50b90a35842dfd60bae49063e3e482b453673d6cdf0cc862a2907ef"
// synthesis attribute INIT_34 of bigblock1 is "256'h04044040ff019574d259dc592abe9b5436bc25676154225435480f552892b2c7"
// synthesis attribute INIT_35 of bigblock1 is "256'h5bd12034800374b8fb72c7ff67f4f74008caee9a68dd2151302caad22611e36d"
// synthesis attribute INIT_36 of bigblock1 is "256'h9002c18543c94934360c6de4670775002618276f0bf1653a7a18c29bf01a8941"
// synthesis attribute INIT_37 of bigblock1 is "256'h93908b662e0ff49d62d480cf7291b4332a1c1ec6212c5035e52258f5000a4480"
// synthesis attribute INIT_38 of bigblock1 is "256'hef3d052e4c8c36e12a5bf0a5eb432cd3bde4635dfe0c372ff689d0dfffc42b6d"
// synthesis attribute INIT_39 of bigblock1 is "256'h031ca59edf36694b9deec570042afced2edaaaab3222423122d26e6b998e7881"
// synthesis attribute INIT_3A of bigblock1 is "256'h4ad85626a2252f9208c2cdae4945815ac55c81f3d0902547fffc002b8114c5c0"
// synthesis attribute INIT_3B of bigblock1 is "256'hf2290fe0e1cb74ec6467c5bcc5a84064aed4b3d524986ea975a0dccf2025d549"
// synthesis attribute INIT_3C of bigblock1 is "256'hab1c227790a3c0a726d5c8e0d07c8ab64a8cb91ae8320ae58197b1f363e6bd30"
// synthesis attribute INIT_3D of bigblock1 is "256'hed47081da1ced33e8e36985ae675908639b6ed12a9ee805df749a41674dba690"
// synthesis attribute INIT_3E of bigblock1 is "256'h1c92319998516b69120de886615e347f74f18465b54e91d5a33fa8aa20f6cd55"
// synthesis attribute INIT_3F of bigblock1 is "256'h429bb01d862d5be1f838800274c7fb722cffb389e997db0826ad4dc98a8d9202"
// synthesis attribute INIT_00 of bigblock2 is "256'h404d518fdf73e8456b301bee20d414886df073095880a620316f4ca125167d0d"
// synthesis attribute INIT_01 of bigblock2 is "256'hf925480a11f071212544ed160948066a1411043bb0944a3258c8226391ff3e54"
// synthesis attribute INIT_02 of bigblock2 is "256'h367d200c5a68fda41e31d4f0c4cd5505125047f11aa2c8072385883a63069f17"
// synthesis attribute INIT_03 of bigblock2 is "256'hcddfe9bc14a7be3bd9f5539c4053dd158b6ce9ba43f68f7839be5429b5951b69"
// synthesis attribute INIT_04 of bigblock2 is "256'h7eed77b6ce4b4c85d434d12953ab4572248b68b08818cd81b329b5cba6d0956d"
// synthesis attribute INIT_05 of bigblock2 is "256'hd36c1b7be3a86b2f55203c469e3433badee6ce8d528b157e64e7e9ec99a5cb1f"
// synthesis attribute INIT_06 of bigblock2 is "256'h8d7db514c82d0ebc0f91ad2aea0b2df44a96098d6717659182815525eaa0bca9"
// synthesis attribute INIT_07 of bigblock2 is "256'h55ae946d5bfdf6a12cb9bd851864babc3aff23211876563e377620b124cd2b4d"
// synthesis attribute INIT_08 of bigblock2 is "256'h9fe9f2d22f79cf9e6152de2c55d38bd55b5a21120979d10219ad098e3bb47169"
// synthesis attribute INIT_09 of bigblock2 is "256'h4b78c208dd0464bb20296615ddd19929800274d3fb72a9ff967b560e4b2faef3"
// synthesis attribute INIT_0A of bigblock2 is "256'hba3e86f46c235991b51f5fa75859fd277f5a394651192ff49b106be0a4a4937b"
// synthesis attribute INIT_0B of bigblock2 is "256'h9d13b2c74a1793c21292c2850680e2af87a9c3a55dfa30089ae1482a0219d51e"
// synthesis attribute INIT_0C of bigblock2 is "256'hf2526cb2b074455ce3eaad363dee1c9a9ee5b03bb492e56d50a6009327b41b75"
// synthesis attribute INIT_0D of bigblock2 is "256'hd0459a6dafb8f2599dbdc5cb98589ce07b2a9e655e386c09002e420019550340"
// synthesis attribute INIT_0E of bigblock2 is "256'h35652af14068648fee4a4b90eeea0c33cddc4b132c213121495075143ba6ba99"
// synthesis attribute INIT_0F of bigblock2 is "256'h5b9590ba32fbe1022a95b492a297e1c077089d1ae06b36965af804c4cebf43dc"
// synthesis attribute INIT_10 of bigblock2 is "256'h994ca740440a1ec89389d5e3fffd23decde16904f5321ec6907f17981e0f1056"
// synthesis attribute INIT_11 of bigblock2 is "256'hc8d2a5c2d1d72c4b9fe7c15aa52a0b20a6250410eb28c285782350fcd47fd118"
// synthesis attribute INIT_12 of bigblock2 is "256'h2fad69afc9a6d096dc79faf718c54ee6fa2fcb79e1e1dee5a3a0233c51cc4a28"
// synthesis attribute INIT_13 of bigblock2 is "256'h7120a430a77f4b9402b2fd09e49b4028cc2c5ee8cd29000274dffb707bffada6"
// synthesis attribute INIT_14 of bigblock2 is "256'hebc54a78125d0185cd09e500c985138c3e08ecdd16adc6777ac9011870f4738b"
// synthesis attribute INIT_15 of bigblock2 is "256'h58b8564363a628084a7546d25852211a2e02b308b810a163ee8269e9c3af05c6"
// synthesis attribute INIT_16 of bigblock2 is "256'h9be6e1db355f2f2b9718000798405e2920a0da82b3d53c48bd2415cccfb31c63"
// synthesis attribute INIT_17 of bigblock2 is "256'ha5c2e750259fa4ad5b0889444798b6d4ba86302a18f32f93a069488a2ab4a7cb"
// synthesis attribute INIT_18 of bigblock2 is "256'h2cc9995d2f46ec55ff96274962b7591b5e375c93b5fe46ba2aa87b9c2cb6b6ef"
// synthesis attribute INIT_19 of bigblock2 is "256'h8dfe66cc22c1404d6151aa2e54dc25a31b6b67efe63eebec1c439328abeccaae"
// synthesis attribute INIT_1A of bigblock2 is "256'h50c62f149c77e174ec81b1cb903404f0da4aa1990c18e617db6811b60c1c8020"
// synthesis attribute INIT_1B of bigblock2 is "256'h71f8256359de3bc663baa97db3b6df7608740a127e34cb84912971d8420ad842"
// synthesis attribute INIT_1C of bigblock2 is "256'h7274fffb297cb6afb5cc985667a57a6e36f0d4e6cc48c858dc6c3f2af1327d0a"
// synthesis attribute INIT_1D of bigblock2 is "256'h8d88b4348b6e807c185175a6f0c9304b0c239ba91c021e4a512851dd0373eb80"
// synthesis attribute INIT_1E of bigblock2 is "256'h496deb3a0aa016275bf7ee55ee5421bfe46d929f74c5c4547a9588dd707f7dc5"
// synthesis attribute INIT_1F of bigblock2 is "256'hbaf314874d5086f4c28306286952391b3cb24058dfd8b30e6e3e3d4d1a7b3bbe"
// synthesis attribute INIT_20 of bigblock2 is "256'h6332c93f509462825cb6f71b29246cabc17507c55800000890eb0092a7b57ce6"
// synthesis attribute INIT_21 of bigblock2 is "256'h5c50121f14384af34b75c3901b7ec4191a9fcd223f4ebd04f8132e32fdac879a"
// synthesis attribute INIT_22 of bigblock2 is "256'h5b1d46fb569b6593ecfd9f4ad4f2a9c66cc822e6de84d86063e259875dfaa548"
// synthesis attribute INIT_23 of bigblock2 is "256'hcc6f44c72187946c71b410838280fd5fb3e250e8d72e25020ab75044050203c2"
// synthesis attribute INIT_24 of bigblock2 is "256'h91bb6610eba91e9a8349f681e00020520200c8888856f3a1541d883aa1b45ac0"
// synthesis attribute INIT_25 of bigblock2 is "256'hdc726da6caf75631c15af5b4c3a708da7e02bf2804be248264d2e0986ba39c16"
// synthesis attribute INIT_26 of bigblock2 is "256'h4d5c038ff2007274fffb951373bddcc833fd9a4d5b3558e45b2882107b7bae60"
// synthesis attribute INIT_27 of bigblock2 is "256'hfa2921a4f523a0d16830876e0871bd6d73a4f4cb604c0d889b9d21221cf8e9e9"
// synthesis attribute INIT_28 of bigblock2 is "256'hf690cf19ed39f09f77fd48699bdd7de0059c5ce763b55ce354ddf8c5d9be8910"
// synthesis attribute INIT_29 of bigblock2 is "256'h012b589a549265246410519b19e56a831ab38074b9a88266c3c1a490dc6d41a4"
// synthesis attribute INIT_2A of bigblock2 is "256'h9dd066071215065c201ebbc9e0ec16f1a54fa3bdc586028e8f3db64c4da14387"
// synthesis attribute INIT_2B of bigblock2 is "256'haf0c79cf6f931fde5a759ebe37fde3ee089dd8de479c8ca1a379f943c5cf6849"
// synthesis attribute INIT_2C of bigblock2 is "256'hb6db9cb80136f214b8ca6e48a13b8d2a3a3c042a3a093e3cd2482e69890cb58b"
// synthesis attribute INIT_2D of bigblock2 is "256'hf48cdf87f39f4e6848ba0808b3c9d169ff79f815ce7708d1b0a4908f2a0754a2"
// synthesis attribute INIT_2E of bigblock2 is "256'ha77471e9e6b7fd7aa13f3690236a86db64d822db00295b1a9a7f68a87bb1941e"
// synthesis attribute INIT_2F of bigblock2 is "256'hece597dceddc472ba84d4b3386586443688a8a1be5acd2fceec699834c12b9f8"
// synthesis attribute INIT_30 of bigblock2 is "256'h1ba24508b12c475b0349f1807274fffb13b9849fd24e90405385e2f1274c6a09"
// synthesis attribute INIT_31 of bigblock2 is "256'h80cce8d6b4581e848d8ef9a294d0dc200a6da861987c6f84c125740d18a33b7a"
// synthesis attribute INIT_32 of bigblock2 is "256'he872e380fd1df29240825a15f567b4951b8d465942d2b34ce87ec99122279320"
// synthesis attribute INIT_33 of bigblock2 is "256'h46acad8ad365054eb4485c7111048726cb7abcbeb7b60e5e273585ecf23ce8aa"
// synthesis attribute INIT_34 of bigblock2 is "256'hbe7acbdaf55898f6e007e95198c0e064b4b8fa18493765bb88f330b2639f5ce4"
// synthesis attribute INIT_35 of bigblock2 is "256'h895835262153b8ed352f7dee26f7cd4431db97131e943b8774f1ac7dbbaa251f"
// synthesis attribute INIT_36 of bigblock2 is "256'hcd67af2ab492d38d2108fc01a5499d8aee49f88502711830660d4f2aaa7eaba7"
// synthesis attribute INIT_37 of bigblock2 is "256'hcb9b68e51664c201ae7c949952dca247e65e46b84f33606b52cbfaaf1857457a"
// synthesis attribute INIT_38 of bigblock2 is "256'h2db59dca041a7b38f2ec5327e06c0640b567ed39609580588aa15544a94a7d56"
// synthesis attribute INIT_39 of bigblock2 is "256'h724ba11781357ccaa14bdb1e3ae191dea2b5ee9b599ccbef7c435d24b61393a9"
// synthesis attribute INIT_3A of bigblock2 is "256'h604c0cc3abbd2b841d28e96845dd0304f7007074fffb58f31200d131896e6196"
// synthesis attribute INIT_3B of bigblock2 is "256'heae853985ef644b380c0754119480c25e0479d08f43092eea0a6a45677a72ca9"
// synthesis attribute INIT_3C of bigblock2 is "256'hb1008bac0e9b3951e8c91e758dade40132f5297029e56233b7d9db6d5cc65504"
// synthesis attribute INIT_3D of bigblock2 is "256'heb8dcdcbde6109a4e16d6add178b110011b714da2b200b4af49878ea1aa6f9e6"
// synthesis attribute INIT_3E of bigblock2 is "256'hcd99e4f5a52fae6c512d1d06719cf554dbea0ec744aab3bfc567f7cfa4f791fd"
// synthesis attribute INIT_3F of bigblock2 is "256'h60cb2eea68f732ecd4df14382dcaa16ea73d48a8618bcc88b5df79e27149022f"
// synthesis attribute INIT_00 of bigblock3 is "256'h91e5346d6d83b51b49298a264720cfe8859ee173d9c0aaf8e879d1ed86fa14f4"
// synthesis attribute INIT_01 of bigblock3 is "256'h0679b003675024ecda2b127e7b4a18cfb0c0a752a15e75a9e022abd4021fbd6d"
// synthesis attribute INIT_02 of bigblock3 is "256'h4b3b9652452c9e9127222f6e76c5285464ba0d68cc18406f0a562d293243c8c9"
// synthesis attribute INIT_03 of bigblock3 is "256'hbc28be9d78657dd1545404e625b1c70698f119ab76c8056749808cb164e1dc0c"
// synthesis attribute INIT_04 of bigblock3 is "256'hb2c044b0d7730bc0c5a09a08451b48292b43dcd10e45000374f6fb72f8ff59f0"
// synthesis attribute INIT_05 of bigblock3 is "256'hcbfb07d1755fb4284bb2db745e023bad55f3e2fdc5eb8be8d8a532a1ee68ac12"
// synthesis attribute INIT_06 of bigblock3 is "256'h13df86502d3fcf298c37fa1d51cfbf3e4508964570660617a1a97fef4153e459"
// synthesis attribute INIT_07 of bigblock3 is "256'ha6aa9c8c8cbc61a52d370f11c1265f0e173c069b36568840e3c3f86ebf445b33"
// synthesis attribute INIT_08 of bigblock3 is "256'h2a44d7f2b4a793e53885e1571453043a2515d8f81a24cb41aefe91602d68283f"
// synthesis attribute INIT_09 of bigblock3 is "256'hafc2af6fde97ad5bc353ca088b273e5efffd168b47522460c6f687bf0dcca9e1"
// synthesis attribute INIT_0A of bigblock3 is "256'h33049bb1d592470480f776bd1aa9912382e962eb2cbe0768c670b86017fb0000"
// synthesis attribute INIT_0B of bigblock3 is "256'h934d11d1279bce99140246c6a3c68983000204511fb974f790445f43cc003776"
// synthesis attribute INIT_0C of bigblock3 is "256'h967f8a3cc2e5b9220f1272aeba5028e58a961a86f42a27603028491110fe613a"
// synthesis attribute INIT_0D of bigblock3 is "256'hfb7232ff4f140665861551fc3d06287f8963c610ae96744854c532e4b9686554"
// synthesis attribute INIT_0E of bigblock3 is "256'h608cee249c0d7248a618df714b98454c8a0ca4bbb82b881edc694d47000374f7"
// synthesis attribute INIT_0F of bigblock3 is "256'h6fff1fa03bd940ef381c18d157c106d55677624be34100816098ff201246d1d5"
// synthesis attribute INIT_10 of bigblock3 is "256'h0162004200001160a644e68880891e9da20fd9f74aecb91b96d965f33d159f5d"
// synthesis attribute INIT_11 of bigblock3 is "256'hcc30a4613065050ebaa1c40b4d7014a854e1854d9791bb8c8942531491194615"
// synthesis attribute INIT_12 of bigblock3 is "256'h25060906cdaa94c1dc8d0352c5c65a118981875c5471677406ac80c419839da3"
// synthesis attribute INIT_13 of bigblock3 is "256'h8cf943d057d339974f9009ea4347cf49604c19db470ee74e2bc0e254c2a906a0"
// synthesis attribute INIT_14 of bigblock3 is "256'hdb849ce2604281820a20df225f550080bf7e9211139aca35efa858db6cb7ec53"
// synthesis attribute INIT_15 of bigblock3 is "256'h6d4168612039431062d783a8b132983a159f8133040900008109800061601b53"
// synthesis attribute INIT_16 of bigblock3 is "256'hdf7b6d2b7eaabb4b9e63def062f08d192eef10fbd857c9e070b7c495501daab5"
// synthesis attribute INIT_17 of bigblock3 is "256'hba40800274f5fb72e6ffadac6e56ad6aa8fc24f41723d767fcdcfbcaa824aed2"
// synthesis attribute INIT_18 of bigblock3 is "256'h8992a1a88129608aed88650a75a0c4a0276c4db5a376690ce4db902c861c5b49"
// synthesis attribute INIT_19 of bigblock3 is "256'he50ea252281d7fd4615f00804596ded669feeec18cfe5f9593dd3a2896db9739"
// synthesis attribute INIT_1A of bigblock3 is "256'h4d4240af59c412072d2545b3976a31a41e4829c000000000990837b58aa4d6ee"
// synthesis attribute INIT_1B of bigblock3 is "256'h6d321399b41842928916cada974840cbd44f1ddd2da9f2c89060f63d6e65116d"
// synthesis attribute INIT_1C of bigblock3 is "256'h3b0390ab0ac8ba197d9f9631f5bc8826d59b5db0cde4a2a054ebb637b89878c0"
// synthesis attribute INIT_1D of bigblock3 is "256'h7d5cf85bb217f8c96abe34408fbc936a659509c36576e73f2f8ea2353bb242c6"
// synthesis attribute INIT_1E of bigblock3 is "256'h7dfeb6fd718ea866318cd0a5eaa748d51bacd0f400c81800f3dfc446d5e944b3"
// synthesis attribute INIT_1F of bigblock3 is "256'h2447f14db95524705e8b242354204088462532804cb04e8834308f1b4d1a1736"
// synthesis attribute INIT_20 of bigblock3 is "256'hcb546ce124ee479d4a25036c32b32ee88a1715a228895248a4d7337aaa397a44"
// synthesis attribute INIT_21 of bigblock3 is "256'hf814234ddc51c760000374fbfb7053ffa0a5b2adad354da8da4606b2c72a305a"
// synthesis attribute INIT_22 of bigblock3 is "256'h54cdd9e53cdb5a9c6cb1412c30982e244a8555a884985b710d8543008904619b"
// synthesis attribute INIT_23 of bigblock3 is "256'hbb61a5718d03444ba7805821eaae4fff0000d28d6e7c0e5eda0997fcb1fde0ec"
// synthesis attribute INIT_24 of bigblock3 is "256'h0aec4cb3907d277aec95cecca1f5122a16c6187287c7000ac122412125db56d6"
// synthesis attribute INIT_25 of bigblock3 is "256'h771b064477d2e23076b2b0936f8b2c1259ce083d0b25aeac8890f6c3e9e2e73d"
// synthesis attribute INIT_26 of bigblock3 is "256'hdd98f43b9ecfa7312dd8aeadd6c8bcab29f5c273b2cbd7dd3dd572e407f7d907"
// synthesis attribute INIT_27 of bigblock3 is "256'hd2427338bd06b64cc8c0807262c8d7ffc802b72353448c2de5606bd7c4f716bc"
// synthesis attribute INIT_28 of bigblock3 is "256'h9a07ce4eedcd708e2531d06069f4f327813afeb0df08faf158785cc62a5cccfc"
// synthesis attribute INIT_29 of bigblock3 is "256'hf2e2327242ff0e9966f3774791c065af663c984bfd5ca4790d3f84d13db5971b"
// synthesis attribute INIT_2A of bigblock3 is "256'h015a020ab8e13e70e2cd2298ff277198f7a84428330ff32b8503b83358045dd8"
// synthesis attribute INIT_2B of bigblock3 is "256'h085005865b4613e11af251e946da036fff807274fffbca12e763367d6278e098"
// synthesis attribute INIT_2C of bigblock3 is "256'h51586f1fa91bc1207916480504b84dbe8a332509249305ade85ca5116847291f"
// synthesis attribute INIT_2D of bigblock3 is "256'h27d5921628e51b39999553593195adaed622d8e729b76eabef593786e5a21f1c"
// synthesis attribute INIT_2E of bigblock3 is "256'h23d7743f825d2ee741679e332c69b5735905e289d2f14cde48016802824c1721"
// synthesis attribute INIT_2F of bigblock3 is "256'h7abbb60d73b468907597fb285f14d6ec1c492c87f053e7e25e30599797ee6f8e"
// synthesis attribute INIT_30 of bigblock3 is "256'ha6058f3c85f3bf73100c52cf422b1277556fe8a4fd0d56c922f6e5fb851fb95d"
// synthesis attribute INIT_31 of bigblock3 is "256'h7742361c2b282d0e5d9386945ab822abc23b2febda84d9f846da4902c73428f0"
// synthesis attribute INIT_32 of bigblock3 is "256'hd07c3242b65859370e143163a25400c2000019803710d018b46d47dc412e622e"
// synthesis attribute INIT_33 of bigblock3 is "256'h39b0719158c91d57b195c6aac9f5cdd1089ad506cfad9dec6844a6bc0f02481d"
// synthesis attribute INIT_34 of bigblock3 is "256'h4ff73514cb5d16a35fccc1b5675767543390f46769315ea2f55627a933256b7f"
// synthesis attribute INIT_35 of bigblock3 is "256'h0cb87146f8d1084b0103db8622e31728392857dc034afd807274fffb7d5adcfe"
// synthesis attribute INIT_36 of bigblock3 is "256'hc752fda38cac62fa861b2ae5241c2a3070758e6599faef7614e134f68f6e40b0"
// synthesis attribute INIT_37 of bigblock3 is "256'h80950187600446296e5c87c5785c3803471b36cca6212ab4b691db9170364d90"
// synthesis attribute INIT_38 of bigblock3 is "256'h3ae3c79ffe2eb9066bc91772420b3e3d636e99a7a325699684878b752d3ea2d7"
// synthesis attribute INIT_39 of bigblock3 is "256'h9f629e2204ee42fa21d675c93c9d6682526fa43b1f049aa0627c95ed2ac3e685"
// synthesis attribute INIT_3A of bigblock3 is "256'h011f3014480098883e3acf2b865fa8577fbb249264b663504f921f565b5fdccc"
// synthesis attribute INIT_3B of bigblock3 is "256'hfd6fe9b21d170224d34990803b306dd4c723a10478015ff411774e832fac2b2c"
// synthesis attribute INIT_3C of bigblock3 is "256'h23463d43abd8c5549307c0bc365ae4f3001b4ea01a20f0473ae3b7284a7a6d21"
// synthesis attribute INIT_3D of bigblock3 is "256'hd5d83e3dee24dcaddb1e2df83d5dd7b7bb78adae913407e9107f90cf9d6b9440"
// synthesis attribute INIT_3E of bigblock3 is "256'hfffb102e25a3e60c141052da95b516dcc81d84e3209cd0a0f617b60f29d56942"
// synthesis attribute INIT_3F of bigblock3 is "256'he81405ade05db1726f443911740e30a2eb7a29832d20e9e844db0304fc807274"
// synthesis attribute INIT_00 of bigblock4 is "256'h6d7148db4002bf403a255b7b86a87e47ea99b0965bc62ee9ded2b5b767be9821"
// synthesis attribute INIT_01 of bigblock4 is "256'h89854a8901440000d000880b824c6b12da9022a72636a61f546e02b8964b7306"
// synthesis attribute INIT_02 of bigblock4 is "256'he3c941e7f14c818c9cf60bccb61e03a8e718d0c7260d5492963372820bd188fb"
// synthesis attribute INIT_03 of bigblock4 is "256'h0fccdca332456122bb79a6504d6587339b897deb7af224ea35bace6961ab3b75"
// synthesis attribute INIT_04 of bigblock4 is "256'h00010268a72fbf77bf151f48a75b27a8e3ee34e0a5a8548370e85fddf9ed614e"
// synthesis attribute INIT_05 of bigblock4 is "256'h1a6406e600103040a806d9a097e2cbc9bbdc4a6ca2286a8529303ae28db7c91c"
// synthesis attribute INIT_06 of bigblock4 is "256'hff3bf27da8b588b28666d6ebbef2d162b2d49d56e9f3fb4db3d08250e2e3375b"
// synthesis attribute INIT_07 of bigblock4 is "256'h696e4c8ba3b2ff53e1c3688340c9f0943ba080ccb7228a6117f3e888ee30ae86"
// synthesis attribute INIT_08 of bigblock4 is "256'h0395fe007074fffbdecd7ad6720040e59de28e866efaeffd6feb3fe3d7cec6f5"
// synthesis attribute INIT_09 of bigblock4 is "256'h4400cb0114919c268a6da06d25166cc63d27844d2465bb6a21225b18498f455b"
// synthesis attribute INIT_0A of bigblock4 is "256'hf937ffc3de50fc03bb332ff38364f9479190b994ab6188c644edb71e9c6d0002"
// synthesis attribute INIT_0B of bigblock4 is "256'h58404943213ca196b9e6624350d4406d78540ebe90013184bbd2f5207bd34d21"
// synthesis attribute INIT_0C of bigblock4 is "256'h74d6ffde48f55b802b6a66eb0df8df6dd48cde6eb46834a0610b78e63a20a6a7"
// synthesis attribute INIT_0D of bigblock4 is "256'h604958a096b7514b237eeb32f1d8153235818dead56c2824bb3ff413b0fe458d"
// synthesis attribute INIT_0E of bigblock4 is "256'hae1a744cff916ec3e1ac81badb7621c8fff8ffffffffffff63ff3f50dea77dd9"
// synthesis attribute INIT_0F of bigblock4 is "256'h5c6b585c75575e7d702202150900e041bf0583b4d8e81c1bf040380881429f1c"
// synthesis attribute INIT_10 of bigblock4 is "256'ha3db8c23cb0d618c72183e31606f2e996bcd725a0de408c79ab04e28d0d48e9b"
// synthesis attribute INIT_11 of bigblock4 is "256'hd37ab98472243797373112d94573cd08784c79626e28971d104e758f0f737a60"
// synthesis attribute INIT_12 of bigblock4 is "256'h701aec5a5a513834000374fcfb7231ff7bfb97f5adfddd4e1277657fadcf84bb"
// synthesis attribute INIT_13 of bigblock4 is "256'hfb400e1c2487a4213dca88116c18ed34ac0d07c08c3d07694c4d0c204d1ba16b"
// synthesis attribute INIT_14 of bigblock4 is "256'h1e1c7b05c3c68321301d7af4ec83c6e381c6e3ee8672080998c8e3e11bffd080"
// synthesis attribute INIT_15 of bigblock4 is "256'he5853b5956c73797196406299781f41bdc0feee93c9acf3a0000b1b640007509"
// synthesis attribute INIT_16 of bigblock4 is "256'hfa819ec5b8356055b2a7630ee9e5324064754a66158ce30435f81217913f8489"
// synthesis attribute INIT_17 of bigblock4 is "256'h2019ca33f22d53629bf768f46a5dd7269affaf4ba836a98388d9c68e723b87f3"
// synthesis attribute INIT_18 of bigblock4 is "256'h2bfbc1442ec6dc6d81b60800195fa8427183bc59d41960d8215858ea8e472a54"
// synthesis attribute INIT_19 of bigblock4 is "256'h8330cbaed1650039ce2a010881eb8fe6176eeb195bb3d8016d319b2988dea131"
// synthesis attribute INIT_1A of bigblock4 is "256'h390626a2106ec8bf3daecba8d8f6a85e79559a237e0f1876cffc59326c90934d"
// synthesis attribute INIT_1B of bigblock4 is "256'h8f3e631c7b32e7554a4c770bb6eb64baa25323b90ef58e20b78b06d71baba26e"
// synthesis attribute INIT_1C of bigblock4 is "256'h831a5315435b6021892c5ab93d41800374fffb72a6fffb57e02bc72a3736820b"
// synthesis attribute INIT_1D of bigblock4 is "256'hd36e204c93016f33d6fd63e869315e2611be148c6d58858d5748e6206f6a4d79"
// synthesis attribute INIT_1E of bigblock4 is "256'h850000803e2896ac9a30679613556b4c88dc8938518cfce56eaa0b296a8d36d6"
// synthesis attribute INIT_1F of bigblock4 is "256'hb3da38aceffaac484c81ccb90ae217d3a203366ad2a505efdc83ea480ba300ce"
// synthesis attribute INIT_20 of bigblock4 is "256'h4663f0216b27d8bad785580fff0d01515e9f0a35bb409467b9f09f3e954cb2ef"
// synthesis attribute INIT_21 of bigblock4 is "256'h0456d13541d182176f460b63ab5a045773dcdeb4ff7196de1b286737f2ccdd72"
// synthesis attribute INIT_22 of bigblock4 is "256'h7e336294172f87b383982bfa19538e504fffe70125ff4831501d0c8f80dba63a"
// synthesis attribute INIT_23 of bigblock4 is "256'h49eec74a62faf452bd31c0b5ea9491870001000400130aae332ff575caec60e2"
// synthesis attribute INIT_24 of bigblock4 is "256'hb3c54ccbda1ad2f989b95cc0e8247bdc38c3796d1a9043d0994fcc4d570ed806"
// synthesis attribute INIT_25 of bigblock4 is "256'h4bd0cc461f7c6baf99cb030bb2e1ce5785460031cea3f86a8209851736fd0544"
// synthesis attribute INIT_26 of bigblock4 is "256'h24a007734c59e62e9a04635b4a20881e5cd1905f800374fffb721cffb1a75167"
// synthesis attribute INIT_27 of bigblock4 is "256'h203cbb48ffe0800b4c693bd05cc1d9119e6169c42040899414946e68820db1a8"
// synthesis attribute INIT_28 of bigblock4 is "256'h0f9f963993d70e55d00047000431432eebe774530ba8e71f7cb094ef5a3d961e"
// synthesis attribute INIT_29 of bigblock4 is "256'h1db7d3485d5fa3b9533ebebd7d5438984d6b4f91b71731ff68f8470484f75ab8"
// synthesis attribute INIT_2A of bigblock4 is "256'he852a530992265e6e7d6c4a122d9d381c1634ef6be6d5c336b873b77e9466cff"
// synthesis attribute INIT_2B of bigblock4 is "256'hc1b0ffffffffffffffff15ff7429e4e48de1d9e91d30b1663fc1f5231ae63b84"
// synthesis attribute INIT_2C of bigblock4 is "256'h5d18d000ea16476294d68b7666c2267c6d22b5b6dd2a176462c1e164224bbfff"
// synthesis attribute INIT_2D of bigblock4 is "256'h4cb6cd8bd074153bee972bb62a68cd1eca3a9c9534ab46c294ee808400510400"
// synthesis attribute INIT_2E of bigblock4 is "256'hb4908c573aea9a64a54d39b98138cc3450f7362c713798d6b1df3dc6ac76f779"
// synthesis attribute INIT_2F of bigblock4 is "256'h6bff242551cb1379b6930eb546c77f822a916be3da1430fabfa38db9d31d8066"
// synthesis attribute INIT_30 of bigblock4 is "256'hed98758db1a0462c176d4d39e5226605835bf81d891cdb498345800374fffb70"
// synthesis attribute INIT_31 of bigblock4 is "256'he8ba1911375b0ec122b8f8b3fd9efffa4002800c935e2d8e1e958483a0051308"
// synthesis attribute INIT_32 of bigblock4 is "256'h0e6281786c1cc7da8b8700468000008ce400b05493fcab6ecd0a45d6511d504b"
// synthesis attribute INIT_33 of bigblock4 is "256'hb91f866bb2e6847b4e117893609e6989341922da809c3ce80046131728106bde"
// synthesis attribute INIT_34 of bigblock4 is "256'haa6d8ad8ba32d772d1ccdcbe180165d3ed4c2e0858eea2d662c6e7792b9fad70"
// synthesis attribute INIT_35 of bigblock4 is "256'hb6db52314680fff0ffffffff6ba7abd836a328ebf738f2214a1884f36aac194c"
// synthesis attribute INIT_36 of bigblock4 is "256'h1a005ff13af79e1527d8c6342bf2867968222a2f4a0c4ca34ecc528c71cf9f01"
// synthesis attribute INIT_37 of bigblock4 is "256'h20bb77a502367a71e5a4a80e131967fadf65b46989c628e73e251c8800006c49"
// synthesis attribute INIT_38 of bigblock4 is "256'ha86ba2e41c1a8145eb5f95879b388ffdb4788b6b25997e65aadd36d8f8f92ff1"
// synthesis attribute INIT_39 of bigblock4 is "256'h034aff807274fffb905da74de5f819f95bfeb0b9a9b9d6ffd2a0edf339559c81"
// synthesis attribute INIT_3A of bigblock4 is "256'h569fee3a99e1a4920d6da08a2d186d466915384d1cc55b661f031788318741db"
// synthesis attribute INIT_3B of bigblock4 is "256'ha06b1a2f8305dab127229f3f4faaf912d987bd9cdb6e28b8100036c221ff4d9d"
// synthesis attribute INIT_3C of bigblock4 is "256'h54ef019bc9e950f632d62a14f8678fc5005d440022002602c330456d0191c33c"
// synthesis attribute INIT_3D of bigblock4 is "256'hedbf743c5ede2bc5329ae8e9475e6f4b3ff28c6f74977b0c851117e3fddca680"
// synthesis attribute INIT_3E of bigblock4 is "256'h8ae85552ecbca15d7ee2ec7ebbb3e52dd9d29ae753f0365fd2bbcb7a9b234c49"
// synthesis attribute INIT_3F of bigblock4 is "256'h7c6d995cb24010c9ffdc15ffa01468f09052e236ce690c51afe891fba98921df"
// synthesis attribute INIT_00 of bigblock5 is "256'h181c0d434000284048088500fb97b0d97ad71dd11ad98fee11cec2caa4a9d682"
// synthesis attribute INIT_01 of bigblock5 is "256'h52cb9ed43ae9f93af69fa028ea1f908c98d1142c69153a10a4773635dc792121"
// synthesis attribute INIT_02 of bigblock5 is "256'h8cf420167499bf4d5838dad41f7a0a74995245fdd623bb9b40ab9e330ad7d769"
// synthesis attribute INIT_03 of bigblock5 is "256'h2f885126415b0354ff807274fffbb9f11c88bf741f5cc84a8d654908e5594e9b"
// synthesis attribute INIT_04 of bigblock5 is "256'hed613bd015fc5ddaeb6c89d8a8920ded288f1cbe6ce62cd1724c18465b6a2663"
// synthesis attribute INIT_05 of bigblock5 is "256'h0a3e3a3d4b67315f20d95f5380921d5034506835f629ee407ba76db7906300de"
// synthesis attribute INIT_06 of bigblock5 is "256'h1d28262d35830d2928178aa1040da51b9ce85100000164120008abc04f50137e"
// synthesis attribute INIT_07 of bigblock5 is "256'hcf4b482057c61c23d4c89a7de2b949978c6c06a3cd67823b1bd1eae4265085b4"
// synthesis attribute INIT_08 of bigblock5 is "256'hc0a7b8db855f737a9042eb14ca2e22b952387bfb5b9d3503e3d507982b05bc93"
// synthesis attribute INIT_09 of bigblock5 is "256'h189a194dbf8b6db682630000fffcffffffffffff7fff2ccdad6a6eaf1b49ac73"
// synthesis attribute INIT_0A of bigblock5 is "256'h8000580000003d337330561b729d963e80bfb4a25c93b2ce779f692084eac3b0"
// synthesis attribute INIT_0B of bigblock5 is "256'h06361146ffa3db841955698d241616363e490dcaab525d636a58daa0c8c21b18"
// synthesis attribute INIT_0C of bigblock5 is "256'h0885e873f84652b15b43349e881d525acf66ae88a9cea6edcf44a127b766c432"
// synthesis attribute INIT_0D of bigblock5 is "256'h24266b6923a3147861ec49db0344ff807274fffba185a8b4a430cec74c700c44"
// synthesis attribute INIT_0E of bigblock5 is "256'h00805a68fd9d7a5d334bd8f4557efeca1ec1a8918d6d209a205e6da6c919720c"
// synthesis attribute INIT_0F of bigblock5 is "256'ha00630a4056796ba7f66a0cdd9283c4ee597283a66bd13ed4f0eae1f36017fff"
// synthesis attribute INIT_10 of bigblock5 is "256'h62803bcf6760da54e91ec8d5830825de016ab53a1418520d1e1847512f86211c"
// synthesis attribute INIT_11 of bigblock5 is "256'h6fea4039a9e7636d07c8e4c1d758d510dfe20162decb297e21120d3d98e5fce5"
// synthesis attribute INIT_12 of bigblock5 is "256'hfffffffffffffffffd3f7aff5b3b886adab7c83d1b97ecae1667b4a4393b6214"
// synthesis attribute INIT_13 of bigblock5 is "256'hcda4a9e8a09e0ab4ed5be5f199cc50b5dbef8542a85b6063db6f4eb62000ffc1"
// synthesis attribute INIT_14 of bigblock5 is "256'h47f562f729a162ff6ab9e99a2359758bf4f1478000053050ae948820338070e3"
// synthesis attribute INIT_15 of bigblock5 is "256'h10c53bbb305abedaabac0ea27d27f769733a247af185a256fbb2fe709331a544"
// synthesis attribute INIT_16 of bigblock5 is "256'hfe65b862df75d58abf9b88dcddba9cc7c674574664a9c832a22d7d00be98a9dc"
// synthesis attribute INIT_17 of bigblock5 is "256'h6d46f507940b24697b6a26a31638512b415b036efe007074fffba03c60af7934"
// synthesis attribute INIT_18 of bigblock5 is "256'ha43907593a04f746fffd02044842c7a7cbf09ee5416994b198340d6da07824b1"
// synthesis attribute INIT_19 of bigblock5 is "256'hd6b8333f07aea00002042aca95d420cc0c20ab1f13a0ebf7bbecb03e504e79d4"
// synthesis attribute INIT_1A of bigblock5 is "256'h5461cd8ac136b38410d5cbb39fc8ae9326b24cefed2c84a1c956bd3a7692693e"
// synthesis attribute INIT_1B of bigblock5 is "256'hb4a1ccd3bc9222f6044ea8131c6955aa6d8296c25aed714261fbc4813e2728e5"
// synthesis attribute INIT_1C of bigblock5 is "256'hc50cf2616ef9e126a4df7a0cd6bfb6614f8fb9b40fedd6bc0bac3f7f57f33d54"
// synthesis attribute INIT_1D of bigblock5 is "256'h09a811523bb889b4152bafa06946371b0021577f07145be1a8e124d18bb136c2"
// synthesis attribute INIT_1E of bigblock5 is "256'h8a89bdace120e9c326dc00c71218848057487ec37f88f0ecd9c0ec36ea11e8e2"
// synthesis attribute INIT_1F of bigblock5 is "256'h0361d4c4e8756647c2325432ab29717ab194e9af0bbae2e3ffa1bc93052d5fac"
// synthesis attribute INIT_20 of bigblock5 is "256'hadff15c39b0651f7bf2a4370feb2d9cd75c74213fad8ffac2f60d37a482affea"
// synthesis attribute INIT_21 of bigblock5 is "256'h6da48d8d5ae0e62c156c0cf1094c6a15e37bc8252b2d5b312a41800374fffb72"
// synthesis attribute INIT_22 of bigblock5 is "256'hf290aa6ae46d189453011a81ae71e3ce12a256d109f04081e2c42c1e88c3611e"
// synthesis attribute INIT_23 of bigblock5 is "256'h5e8e38230640a00080a414e9ad74b333465cd907747c27c9d3948dfa91a2c242"
// synthesis attribute INIT_24 of bigblock5 is "256'hde3e7cd3841645ad939f352910db3bca115673f356e795a90be99a56a8744553"
// synthesis attribute INIT_25 of bigblock5 is "256'h0639aa9098faf88b4b50cc1b6c8d07e76cca6b7cf80efeb00c172711de3e7299"
// synthesis attribute INIT_26 of bigblock5 is "256'h5fc0f6a18c70021545c3d55b0233a1685b8a127d72e8a9c72d37d5aaca2bdd2e"
// synthesis attribute INIT_27 of bigblock5 is "256'h654cf0ed4389457fca3ffc0f225805d04ee639f09bcde265660757a238db104e"
// synthesis attribute INIT_28 of bigblock5 is "256'h8ca960b1298ed1560f37c3b9cc54b5a75c1a23cc0b681ba802dd300000251478"
// synthesis attribute INIT_29 of bigblock5 is "256'h067e28c4e55b588a5fe894cf7b15905d11e5611ebd08559e26e2ad80f6697b4c"
// synthesis attribute INIT_2A of bigblock5 is "256'h800374fffb72bbfffe55165398dad2ad6b98a18890743b63f1c71746ce0df911"
// synthesis attribute INIT_2B of bigblock5 is "256'h8b7238d113086ddc7a8d1460262de16f0c6846767720237bf822884ddbb9c060"
// synthesis attribute INIT_2C of bigblock5 is "256'h39df2f7adec5e69988855187e5a557a6e38d2d2824000e48d887e15abbfce774"
// synthesis attribute INIT_2D of bigblock5 is "256'h734cb2ad3c35bdba4602000004109490c4658711d5b8d8d32db0d81dff2528a4"
// synthesis attribute INIT_2E of bigblock5 is "256'hbcbf96e19ebe9453449957144b50f1b792573462183e72ea5ee46d8363d64271"
// synthesis attribute INIT_2F of bigblock5 is "256'hbdfd3a9aded572cab4e3caadfe5e65e71b88fa15b24db49776a6d0607d7f1a47"
// synthesis attribute INIT_30 of bigblock5 is "256'h52c80a2f6590a3cae46d1024c76e7aed3a1bf5fbb8d30a2d9fff53e63d91c28b"
// synthesis attribute INIT_31 of bigblock5 is "256'ha3b397c4000285a048028217c5f8bc14a5d858bee21713ca5d4ab46528733991"
// synthesis attribute INIT_32 of bigblock5 is "256'h6a7b75d1b4a975a583cddad31377ef8b54d96447066b87bb2ba5d37ac158224d"
// synthesis attribute INIT_33 of bigblock5 is "256'hbd3198bf1f1c0cc1ef18b62800e4d07c6ebbe68232785819a3e94614d67d73b1"
// synthesis attribute INIT_34 of bigblock5 is "256'heb2c5b394a49800374fcfb721dffe9ebf30ed6d924f863017a43d8abd1f06261"
// synthesis attribute INIT_35 of bigblock5 is "256'h52461623abd4d0e5a9db93096da8998defe047a4136d0ca12326670d636b7821"
// synthesis attribute INIT_36 of bigblock5 is "256'h9b0a008a16355fb12a01f2a130a3efae4f4d1e13f44ead625247c2cbe1dddb9c"
// synthesis attribute INIT_37 of bigblock5 is "256'h214a57b64912c595b05a7d35613c5b980b15784f0d61f4e9073142209b2cd077"
// synthesis attribute INIT_38 of bigblock5 is "256'h06e5803c56c988267826c75450faf95bc38e5d503c64efb09b88ae5857954d5a"
// synthesis attribute INIT_39 of bigblock5 is "256'h50066f9f47df650f0ad557731993d2b64ea9cdfa952330f1de6d2d4788f2675b"
// synthesis attribute INIT_3A of bigblock5 is "256'h196560899c8077b46db8832420004f0828bfbfdb676512b5073748e923e53fdb"
// synthesis attribute INIT_3B of bigblock5 is "256'h049c00405e08d1a5aa17c872b63205588172b93a1f21ada87cd43c26d6884e49"
// synthesis attribute INIT_3C of bigblock5 is "256'h641ee0c39de3af2c0950658dc5970d3b2884076e37ac291f194c7370c65a9252"
// synthesis attribute INIT_3D of bigblock5 is "256'h52ddda1f32ca2a4d72752ea29ed51111f6ab141159908e1799331858535910b1"
// synthesis attribute INIT_3E of bigblock5 is "256'h570042bbc822e95bdad11b44800374fcfb7032ffe5fce3df3f6db6cf5e6b115c"
// synthesis attribute INIT_3F of bigblock5 is "256'h5c6d71b7012400006b08e8f41d7ff8fdb4a06d5c9c8cbae04620136b4c49c70e"
// synthesis attribute INIT_00 of bigblock6 is "256'h00a179579a672a3a3c8b064989c3b566b2c8ec4ad1c948466d544176451ad07d"
// synthesis attribute INIT_01 of bigblock6 is "256'hb0b70913545078b91a903d78b22a97c1a40d79a25dd8c3028b2aa609a474000f"
// synthesis attribute INIT_02 of bigblock6 is "256'hff6e3d2896cd1f9dcf843b6743fd51a96ad3d841393b3d39d3f9c9d1dc650633"
// synthesis attribute INIT_03 of bigblock6 is "256'hf6c16044c94fefa11d8a1c728d55cdc8cd4d302ae9979249f67745a2ba06436a"
// synthesis attribute INIT_04 of bigblock6 is "256'h0a85dcacf1ea3dc63abdb0483576a492a000fffcffffffffd7ff4725cdfff7e0"
// synthesis attribute INIT_05 of bigblock6 is "256'h46e8de4c1b9b9b5b0123704083408d1650c6ee269dca02a707f287ba8c5920f8"
// synthesis attribute INIT_06 of bigblock6 is "256'hadf65ded6683910567e5f987206f0cb13bc590e6e5dcdd17697693fda4d0e174"
// synthesis attribute INIT_07 of bigblock6 is "256'hfbdd3810c865ea54952c0b3003e5b5fe4e8beef9a228f6f2c3ff79c0494b7bd3"
// synthesis attribute INIT_08 of bigblock6 is "256'h66e70905820b25077b3a29c31d68b1eb45590370ff807274fffb7ca3d35a224f"
// synthesis attribute INIT_09 of bigblock6 is "256'h1d1e07d03cc4e743238d2019e900352cfed6d9db75ab1c38e8060dec809cb0e7"
// synthesis attribute INIT_0A of bigblock6 is "256'h2a0712e91283000055003ae377540082f6cd1416836f62b6f8d3b0865b3a73d7"
// synthesis attribute INIT_0B of bigblock6 is "256'h347d1a5d333249149d3b3a58abafa7093d98ddb22e9c2a58771d11ebd9fac392"
// synthesis attribute INIT_0C of bigblock6 is "256'h1fc5dc3042e0d8296b32c54592e919861501f6f033f3bd59c5eecb58a94b3773"
// synthesis attribute INIT_0D of bigblock6 is "256'hbfff55aaddfd0d338df77ec009eebee61d90f71f5ca2bcd4683cfbdc036a7dc2"
// synthesis attribute INIT_0E of bigblock6 is "256'hc748477fff49e70a0da5bfea37388eda116d384aa0737241c6ca5491fff0ffff"
// synthesis attribute INIT_0F of bigblock6 is "256'h0ec1ce84a95237098ba382dd7155c782580f9707d01d0003b800c61e592e34ee"
// synthesis attribute INIT_10 of bigblock6 is "256'h92580619ca8b1dd721c834696981a67829eec54ce40496954860c9bcd1e63c70"
// synthesis attribute INIT_11 of bigblock6 is "256'hd002483d1ad8b68f0c34967926181735ec726579ff32c7192c919116116b3bbb"
// synthesis attribute INIT_12 of bigblock6 is "256'h0d6c4090a4b366e77d03284b0d855b3725631798b1884d59037eff007274fffb"
// synthesis attribute INIT_13 of bigblock6 is "256'hf51ea8e88421964aadc9ad0a1feec7a0c3259492f230b38ed3d658680969dc93"
// synthesis attribute INIT_14 of bigblock6 is "256'h99b2a562c440ab84721e57250000e500fc1c5cc485a64f9f2f18d51842e64385"
// synthesis attribute INIT_15 of bigblock6 is "256'h7d195b265ea59fdc9018adfd5b48168412ef1d225160066a96c63dbd95720e8e"
// synthesis attribute INIT_16 of bigblock6 is "256'h83246103dec09e45013e83413e8d67309950d5228eb33219e2fc4c5e7103bc82"
// synthesis attribute INIT_17 of bigblock6 is "256'ha6da0bfff8405fffcf434d3a5a1733c3e921545ca93d237381ba2f7c63dd0569"
// synthesis attribute INIT_18 of bigblock6 is "256'h412038680e65b81a48527b5bd8964e1b1deeda43810d0485212c0aa4f10e0924"
// synthesis attribute INIT_19 of bigblock6 is "256'h75ca3b6b4a8bce0f8ec2c762750c0aacae154e5660f3c3c5426124032aad0000"
// synthesis attribute INIT_1A of bigblock6 is "256'h50ae976305cc4d99fe1a39206f7609cbb9f7fa202f97136f9c4e8286e4b5a58e"
// synthesis attribute INIT_1B of bigblock6 is "256'hff807274fffb34cdd42eb0e26182801092119d0024efb61e58972f763235b4b4"
// synthesis attribute INIT_1C of bigblock6 is "256'h3ccb8ca1c8340d6c607d20756666e4e3064c05063b3323231f98998845590364"
// synthesis attribute INIT_1D of bigblock6 is "256'hf35e124ba345e27131abea472e4c1a038b9cb3ccb612fdd1c105baa05a93350c"
// synthesis attribute INIT_1E of bigblock6 is "256'hc75a3b1538d9adadce66cca4b76b1b4a2b4200000060cc0a333f34a935bf687c"
// synthesis attribute INIT_1F of bigblock6 is "256'hbd965b5d408713428cd51b54c86edb84c7954eb85cdbb9a39ead1c3a09dc9ea8"
// synthesis attribute INIT_20 of bigblock6 is "256'hbd5b10bde77b79430bf835ad2799c7b13339087a8ab8534033bf9e322efe3fe5"
// synthesis attribute INIT_21 of bigblock6 is "256'hfffeffffffffffffffff5257266032029d2cd8298b4a3a69901ebe6a14b2dfcd"
// synthesis attribute INIT_22 of bigblock6 is "256'h0ee58b60002a6000d20473d4d73841d117db4b8cb6014446a89a1da8bc98ebee"
// synthesis attribute INIT_23 of bigblock6 is "256'h49665cf27138f232d6a2792186c8c0de02b16b1d25e6db9abd6fca738e712a79"
// synthesis attribute INIT_24 of bigblock6 is "256'h7b77df585b3b6ea3b4fca3133e89536d28d71ccc2c3189dd13dce289cbacbc42"
// synthesis attribute INIT_25 of bigblock6 is "256'h99e93d58034dff807074fffbf7c3f23e7e79bdffa57efc7d1ddf29ff67cf72fd"
// synthesis attribute INIT_26 of bigblock6 is "256'h80683d8960f0a740986158640a6ce0921876626644e3580c2cc27b1624c31bf8"
// synthesis attribute INIT_27 of bigblock6 is "256'hf035db04af5ed87f96fad0f9ebc1be6aaaab25ea16ca7d41f0343ff023ee8c59"
// synthesis attribute INIT_28 of bigblock6 is "256'ha905c998ac6c9104819349d04152dccda93338049a5083c9005200002cad7e05"
// synthesis attribute INIT_29 of bigblock6 is "256'ha25e0d4b258ea865bd474eb1863863a6a09188921703e10fa26e0a84e47a844a"
// synthesis attribute INIT_2A of bigblock6 is "256'hec87cf15b3e8c1645eb66a99e1a71990927520af5ab6772319640ccf140c75aa"
// synthesis attribute INIT_2B of bigblock6 is "256'hdfe78d6a4ff78fbf47ffd69f8861dc55345e9a1da56756efeea2891d4cd3e32a"
// synthesis attribute INIT_2C of bigblock6 is "256'hfffff03f18a3f838fd40d4fe29554819ba085ae4410a051b325ad072e719aa14"
// synthesis attribute INIT_2D of bigblock6 is "256'h45a300fb010d6698fce042489f0e423474a44d857a14892990910e6a2c4eff67"
// synthesis attribute INIT_2E of bigblock6 is "256'hf354a1aac5717ad87a3ac7e55abe677648660e0f7df6b094139769961368b2ea"
// synthesis attribute INIT_2F of bigblock6 is "256'h121941fb2817e61e58b9ae4b800374fffb72b7ff0883da169026705a393280e2"
// synthesis attribute INIT_30 of bigblock6 is "256'hc98034b4a2e7be801f466b4b2c0a00c69860ec4a5d078020f4f40d620e39e920"
// synthesis attribute INIT_31 of bigblock6 is "256'h5d9c293429d61d67b0adfc9f154509ee8e98902e03a10fd67b538729872e11e0"
// synthesis attribute INIT_32 of bigblock6 is "256'h58fd212800c909b54609f1688bf3485c470575bdcb0a6f333fa4168d887aaf53"
// synthesis attribute INIT_33 of bigblock6 is "256'h9f371a8c574e86ab7a28a6d555cb4356b98c8a407834a449741010c2624598c0"
// synthesis attribute INIT_34 of bigblock6 is "256'habd265b672925ea5131d84478fc988c9f61a4edc8245132b538ed0cfb11b8384"
// synthesis attribute INIT_35 of bigblock6 is "256'h0b9fb70e7cf1d7a3bcec235a7543642ec8e5c6c11adf9ad97546dd3cda18bed7"
// synthesis attribute INIT_36 of bigblock6 is "256'h4359fec2ffffe07f0c176eea21ca3063ec2ce7ffccbe76e60fa696d7f9d864ff"
// synthesis attribute INIT_37 of bigblock6 is "256'h13b439ce58911a5552e75d224d56d65ca5c10e486ccb46905cd0550aab228f47"
// synthesis attribute INIT_38 of bigblock6 is "256'hd4750014ee567ea6bd0e7c58d4db550d00f2cc23595b2a9f472b7bbe23c8fc42"
// synthesis attribute INIT_39 of bigblock6 is "256'h915a1abdb000d2c703ca004261e05696c43f800474fffb72b4ffa6105c07dd8b"
// synthesis attribute INIT_3A of bigblock6 is "256'h15524e72a1001160894e684c974638ebab5c7cc500f31ef02b4b0e8f800119a7"
// synthesis attribute INIT_3B of bigblock6 is "256'hf3d53a3b207ba91a6beeffe1dcf9e16a8ec5683ebb7b97a9aa5708cd758d212b"
// synthesis attribute INIT_3C of bigblock6 is "256'h39cff7dcb7a4394f7becdf3e13b5a99f801cab765414f1f25f2d36cdc543d455"
// synthesis attribute INIT_3D of bigblock6 is "256'hf30a10094744cb765dd8579452b91a0eefed7f95b6db1a8d0138400116c1ea83"
// synthesis attribute INIT_3E of bigblock6 is "256'h48653913cac38c413a850ae70c40955a4e97226636f5b205493414bd62ec4b59"
// synthesis attribute INIT_3F of bigblock6 is "256'hc9ed3189436bf3ae237dd82893820ed84c9df6120e360172fd31bcbfbeb25f0b"
// synthesis attribute INIT_00 of bigblock7 is "256'h50bfa06d61cedd95db5372a3acc54815de7a9455ef212c6534653bddecd3231a"
// synthesis attribute INIT_01 of bigblock7 is "256'he3444672c7ddcab29cc9daaef576a349bac1264d34bfe36dd904740657eb5bfd"
// synthesis attribute INIT_02 of bigblock7 is "256'h2914f88bd4b88a49419351c48c2257564e38fa6f93726c4797a64824eeeb252e"
// synthesis attribute INIT_03 of bigblock7 is "256'h690d4bc8a3244b794c2d9400cde2e2fb0a1e3100de67243c80037490fb72c1ff"
// synthesis attribute INIT_04 of bigblock7 is "256'hfba5747f2afe8fd8e08916657a5d987ba3ac18731ab7f8914b23a8941119ef28"
// synthesis attribute INIT_05 of bigblock7 is "256'hc66f3c5e906f54dce1acdbabca6e7cf7476dce27e34959c7c762c3f9a59ff447"
// synthesis attribute INIT_06 of bigblock7 is "256'h5d50d147a7d3abbfb55a16629c042bf8b692d3cd4356800371cdfdd0bd1492bf"
// synthesis attribute INIT_07 of bigblock7 is "256'haaea77d6a46f100b9e54cec7447c32ba5a53038792e8d883e44f6646e47d8ac4"
// synthesis attribute INIT_08 of bigblock7 is "256'hd11e32eda4bb4da23d7f6fdd87508ee6a0d8558881e31116eb1865fbc4c9fb04"
// synthesis attribute INIT_09 of bigblock7 is "256'h75552dc2f13affad6a7954dc9137b0987cc5ecd6b2a97d1aa6652dde90f486ba"
// synthesis attribute INIT_0A of bigblock7 is "256'h4c894b098837f848ba198c0cbac555ec1a94a9d74917e6dbac5a20b445002e85"
// synthesis attribute INIT_0B of bigblock7 is "256'ha8ae266153c66f6a3a5623b9fc0d35772f0f4219a0cfc79009a20027b700526d"
// synthesis attribute INIT_0C of bigblock7 is "256'h749cfb70cbff354ae58bea0f81365d54fc390e4814fb7bb5b444b19e7d29e87b"
// synthesis attribute INIT_0D of bigblock7 is "256'h60480088efb46b0d5408a5bc277d0bf52732ed00837bda1be91b5f69293d0003"
// synthesis attribute INIT_0E of bigblock7 is "256'h2b594b8f6acb1fec41c21496f075a4ecbbbd4e7c7ef25afc641fa6d41d5ebffd"
// synthesis attribute INIT_0F of bigblock7 is "256'h4e81a1930afe396354ec0ab478c1cf7a08a8494ad3f46da5c91b158121e29d91"
// synthesis attribute INIT_10 of bigblock7 is "256'h0e08bce20f5d476c79d1267a63fac8bfbc8fe5ea0da1a82040204e3604c94b64"
// synthesis attribute INIT_11 of bigblock7 is "256'h353a675aa36f78154478d83add1f30a757d84c3f8aea6b71a246d7afbfc72d1b"
// synthesis attribute INIT_12 of bigblock7 is "256'h0965cc43810bbbaf4b42fecfcecc992e2621e7d19bd01915209d377ddff83b11"
// synthesis attribute INIT_13 of bigblock7 is "256'hd908e2690022930a86acbd5d2032b4f849d2c89c6cfd38364bb9b6db0f314019"
// synthesis attribute INIT_14 of bigblock7 is "256'h4ca9d7f85acb8078224bc5b3d433eb5faaa7099594530d8091b894eda9b4053b"
// synthesis attribute INIT_15 of bigblock7 is "256'hb9276dd06795fd89743727597d34374007d1eafab2903f8a792ff99f93873309"
// synthesis attribute INIT_16 of bigblock7 is "256'he9892edd030ba9007274fffbed6f57dff3e62c76453696efa51d53f7c8a514be"
// synthesis attribute INIT_17 of bigblock7 is "256'hcf004b9d9b606e8709c0e8200deea867945877a4e957340b04657bba1da32d9a"
// synthesis attribute INIT_18 of bigblock7 is "256'h9469c79491e0c20d77d557d0e0c62d4a22769b68535bb06eb4ee1b6d09470751"
// synthesis attribute INIT_19 of bigblock7 is "256'h9cf98e439755c3d21c972d3b2a45c2b238f427bae7ad2b97dad99d6580043916"
// synthesis attribute INIT_1A of bigblock7 is "256'hbca913beed12afe536abb66198870856757ece94260c75f32827c895b514f4a4"
// synthesis attribute INIT_1B of bigblock7 is "256'h9d281cd915a177ba7f1322b7723ca683c31c5d21ca137f4cb9554cfc4ff9c304"
// synthesis attribute INIT_1C of bigblock7 is "256'h044b4748fb7d03820ebbbbd4cf57e964ee289703662701536d2cd91b4a856124"
// synthesis attribute INIT_1D of bigblock7 is "256'h2c75b91871e6f29f96bb94fa071dfe8fdbb65fb8495fa0b74358288840008512"
// synthesis attribute INIT_1E of bigblock7 is "256'heaccd43d19fe6d992318568a038b5756c50287cd43312b71756e3805f9883814"
// synthesis attribute INIT_1F of bigblock7 is "256'h4e46a611008928f0b03524f9d86f5ac60b920bbde516d2e57746cff9e9e8decb"
// synthesis attribute INIT_20 of bigblock7 is "256'h7bcd1e232afa68cc4d5e0308b8007274fffb55cae85f08c56b0471183ce2db51"
// synthesis attribute INIT_21 of bigblock7 is "256'h954254baf3c648e08ffbb7d1de918e1834128defa875087a79a6512f020c0022"
// synthesis attribute INIT_22 of bigblock7 is "256'hadcf2c90040853317dc35247b66d47342e7b7b94acc66ca732bed1b646890025"
// synthesis attribute INIT_23 of bigblock7 is "256'hac588a234655e22eee9ba09747735343a4610c7ae5ea9a28345df1e9145ce5ab"
// synthesis attribute INIT_24 of bigblock7 is "256'h969036d7d99231220022e04cd274e1775352c8bfa2c2ef1ea09af96dace8046c"
// synthesis attribute INIT_25 of bigblock7 is "256'hba844008adb410e3892082b11ab5f1c4e9ac7ee5db12c72186f00103613da149"
// synthesis attribute INIT_26 of bigblock7 is "256'hc3068acae0c50afa1c018f6deb5de5faa4b8b40cc5c76d29cea56f7d16554cd5"
// synthesis attribute INIT_27 of bigblock7 is "256'he09ff5af19c8bd969105c5b32b34a79788c7f19a71fc07eea1c00eeff88de960"
// synthesis attribute INIT_28 of bigblock7 is "256'h159babd691b494dc9c2d40066e3b9fd89de1bf7a87eaeadb40d205f8ee76eb6b"
// synthesis attribute INIT_29 of bigblock7 is "256'h0e1b84e1002692244f48c60bc7065c63e3f8465cfe18e83a706e3d3e8c9257d7"
// synthesis attribute INIT_2A of bigblock7 is "256'h38df020b00237b9d1e833d38e9e541dc02e4c3807274fffbe4d6563ed6226c9b"
// synthesis attribute INIT_2B of bigblock7 is "256'h684d4b3aa28cbb5a6ce4a4931a24211b50d3cd9109a074530c6e6085acb67344"
// synthesis attribute INIT_2C of bigblock7 is "256'h7d9b3fc6727a97fc11d265cbe40b50d60fb63302931b62a8218fd9da543ee55c"
// synthesis attribute INIT_2D of bigblock7 is "256'h6b5948db1a6528bbe208154d76c613a8f04f9f0eceba7418caf6e84d6fdcf3fe"
// synthesis attribute INIT_2E of bigblock7 is "256'hd1ac0005c022505d2e1bb07cccfca31fa0b6f21ce906b210b711080c52ebacac"
// synthesis attribute INIT_2F of bigblock7 is "256'h4ca70a6cde388407125c181d0c7f334a54475d614c9359da7b16667b54b91ba1"
// synthesis attribute INIT_30 of bigblock7 is "256'hee93dd947f9c4a4caa8b5a8c7a6a9e2a744bea3502ebddc4a15daefcaea011ca"
// synthesis attribute INIT_31 of bigblock7 is "256'ha36d9032e008d9bb6fb8fe79f12039334366dd0d5350a221e8b735ec771fc81c"
// synthesis attribute INIT_32 of bigblock7 is "256'h20805f401600b6ee964379ba10a2382089401706456298ce4c0f027fe67db4dc"
// synthesis attribute INIT_33 of bigblock7 is "256'hc5bd990f31efbb8ddd782da015323cdf88d675ffdd81bee10b3fd4affbcc0aa0"
// synthesis attribute INIT_34 of bigblock7 is "256'h2884a4af75a7d93d1e4b00c5bbad1fc2126a692c49dd02ebd3807274fffb3839"
// synthesis attribute INIT_35 of bigblock7 is "256'h92d9d35cafe5179a1e116a1f63397f73a244c4e43abe2539ae970990b4738dee"
// synthesis attribute INIT_36 of bigblock7 is "256'hcb76184b037e87e343bf27f57879a1baf5d29f4ee5e54cab893be3fa65b3d232"
// synthesis attribute INIT_37 of bigblock7 is "256'h457584d600000024ea00449f83afe6d40758f5708e0947ee2492538922244001"
// synthesis attribute INIT_38 of bigblock7 is "256'he2a29a46459bcaa941c6496407032b97a2a19835b8b97c7eaf50ac6c652789e3"
// synthesis attribute INIT_39 of bigblock7 is "256'h2a397b8f6fad51dc20e4f5e6dfb5b79aa76908a8c7e2ac66cf765a850eeff4c4"
// synthesis attribute INIT_3A of bigblock7 is "256'hbb96f47797d30d980d8db5afb1b157e2ef6b824fd9ce97d65769f7dc6792b3e3"
// synthesis attribute INIT_3B of bigblock7 is "256'h0091a5801f9004c1d0f41c3549c5ca8120c46a772492405106f8b149d5fbf45f"
// synthesis attribute INIT_3C of bigblock7 is "256'h697e45558abd54bcb6ef35bf79fc1442203db1ebe8565c85180b8063202c0000"
// synthesis attribute INIT_3D of bigblock7 is "256'h7074fffb4af54aa26d771bc11d3f5c46f47cc1f2590944dd7eefefc01388cdf0"
// synthesis attribute INIT_3E of bigblock7 is "256'h9879f411076de85a20726f46353b0a0c00c27b7a20833c5ad1854bdb0313e000"
// synthesis attribute INIT_3F of bigblock7 is "256'h2100ed05e66aeb22a7978184c06879b191799f91e267d5cdacf649bb72b9b78a"
// synthesis attribute INIT_00 of bigblock8 is "256'h7de83a5f3ba1735d0572cc4dca3b1581d5f5040f580060554c79c55d1380e466"
// synthesis attribute INIT_01 of bigblock8 is "256'hef8c22345ee95a32cd4261f435bb5a39f1daf7be942eee9074dc00060800453a"
// synthesis attribute INIT_02 of bigblock8 is "256'h331cf2762dcd31f23f0c32b78c67d57684a8bd3112079ce442446ff4c322b644"
// synthesis attribute INIT_03 of bigblock8 is "256'hb223867b244dde2d82e53e51986d401600d4edc56d0de4bcf8df864b78f0ff99"
// synthesis attribute INIT_04 of bigblock8 is "256'hb02b339e3e8405cf4ec6945a567bdfddffffffff368deddcd2fff4775edd9fab"
// synthesis attribute INIT_05 of bigblock8 is "256'hbbe2e1431beb1f54faf422605632b9200cc1a5f10b8a0d2d0000f68062c3422b"
// synthesis attribute INIT_06 of bigblock8 is "256'h136aa80d0216385ff8280963907e16eb69c2ee421f3a265653d8a05c500e0867"
// synthesis attribute INIT_07 of bigblock8 is "256'hd949854e000374edfb72a5ffcf3223531ebde67b18a61eecccbd411cdc540330"
// synthesis attribute INIT_08 of bigblock8 is "256'h5329aec30dff700a3324aca45d877720262033654d2d46482718a1cb4a15e933"
// synthesis attribute INIT_09 of bigblock8 is "256'h753ac1c6558a108b1f763fd5d34a51b6512805ab2a9865d1f4ff4cede211fc0d"
// synthesis attribute INIT_0A of bigblock8 is "256'h08a75d468ac9a68451fbb39e4ccf386da0532e2ae95600300000589c26092505"
// synthesis attribute INIT_0B of bigblock8 is "256'hcfddacd165e5c46d1fbfacfda376bbcb2a01befe3647b16a004a5b59ca716cc6"
// synthesis attribute INIT_0C of bigblock8 is "256'hfff3b55f24dfdef3fe6228dc997fbe67bebe5944ff1578313cf0a7f95dbbfc83"
// synthesis attribute INIT_0D of bigblock8 is "256'h8206ffff038454abd6bfe4eb11ff4563242d1d2d2e73fcabfb4f77c717a7bbe6"
// synthesis attribute INIT_0E of bigblock8 is "256'h4d6218d60000010007b4f7619038536b2694a3f24c7e6342d0051059b4a7e24d"
// synthesis attribute INIT_0F of bigblock8 is "256'hfe00d9d8724af227025ba9bdd6b4309f3e9723c327159f0c3ce39cc09f36a2a1"
// synthesis attribute INIT_10 of bigblock8 is "256'h12a2d88eca10bbb98ade7ce23cded69d2c66b54b0fb8c52f9330dfad9b467cbd"
// synthesis attribute INIT_11 of bigblock8 is "256'h21db5a15e933d8b17134800374f4fb72acff973f7befd14a0d4fa5a3ed721425"
// synthesis attribute INIT_12 of bigblock8 is "256'hfd418d62baed55e0e64ed47f295c260cec4c57066d2866240d624cd926601224"
// synthesis attribute INIT_13 of bigblock8 is "256'h264120f1b66b36b5ce2c42fa3b683a1699ea3460dac8693464638346b325c182"
// synthesis attribute INIT_14 of bigblock8 is "256'ha4ab8c02ad9ccf581d4965195fadbb3e3b2dec6b47a98474f340a82f00500000"
// synthesis attribute INIT_15 of bigblock8 is "256'h76179eca1d6df64adccbb64effb78e8baca54de94b6aa3e73da4e4076ecb2b4f"
// synthesis attribute INIT_16 of bigblock8 is "256'hfd6f141be7c6e7dee7e998ebd1488b512b99e52618b106350dc375a478e0552b"
// synthesis attribute INIT_17 of bigblock8 is "256'hc7a79859d1962d24fedcffff55ff49ddd5cbc32bff1e0db439ac0cbebcf5afc0"
// synthesis attribute INIT_18 of bigblock8 is "256'hcb4201649e9a5ee07a7d1fa500060000106bc595bf4f06ad0fd4914a93796aa5"
// synthesis attribute INIT_19 of bigblock8 is "256'h138ff573611c9e80d61d33868c2a66b29c755e12480c86b3e8a02351c8e74ccc"
// synthesis attribute INIT_1A of bigblock8 is "256'hb4474a21ec99079a3e9dd073a665129ad1711765dfc96e0f9c95d2ae60772a63"
// synthesis attribute INIT_1B of bigblock8 is "256'h0d718634f719a1ea4a19ec34d799c14c800374fffb727cffbb1e9d63998bc72c"
// synthesis attribute INIT_1C of bigblock8 is "256'h7d296e8f2a71ae144744d62841e44548f168e1b766186bcc63076fe0e7b0275e"
// synthesis attribute INIT_1D of bigblock8 is "256'hf48255f10000e700a2946e52834e936258901c8bfa94a336fe2bcbc25636d757"
// synthesis attribute INIT_1E of bigblock8 is "256'h4f96a4aec4c6bb7a33577b10a2f25fc3ae38c71e547b886c813ea78c1ef17470"
// synthesis attribute INIT_1F of bigblock8 is "256'h1826db3c41e519b0ae82d2d4bcbfc42eb4a5c76ad670cf651233618749fb5b3d"
// synthesis attribute INIT_20 of bigblock8 is "256'hb1fa20084741b2493fcb98a4357b3223dd2dbc8e10904e392745b9c11ac65cc5"
// synthesis attribute INIT_21 of bigblock8 is "256'he303152c88e0e0eb1891921c8c90fa8cfaafffffffffbfffa4069ef740c56ce7"
// synthesis attribute INIT_22 of bigblock8 is "256'h313a710d8b483561461678a972714de68edaa0e902b2000026201fb84ca52d71"
// synthesis attribute INIT_23 of bigblock8 is "256'h15b14c7d309231c48504b06914473c5abc535e42715499425613c22ce2218045"
// synthesis attribute INIT_24 of bigblock8 is "256'h15f1e3290a993fabe5e794c5d9353a4cd252d8d0e56c5e116b77b5398accf3cb"
// synthesis attribute INIT_25 of bigblock8 is "256'h752067a40b5c4d798918e31981dafa19ec1b5719b74d800374fffb701aff142e"
// synthesis attribute INIT_26 of bigblock8 is "256'h888d8607bbf9866ef30a08567195b9ac8924216e39f2bd51094097a56b886387"
// synthesis attribute INIT_27 of bigblock8 is "256'h44da816e6609da1c7b0700014300988db9e7e0a915f015939e8df38aa0a81d3a"
// synthesis attribute INIT_28 of bigblock8 is "256'h77c73e1b3b424089636c478535051813d9965f745d80230c1a347cc7f4c031fc"
// synthesis attribute INIT_29 of bigblock8 is "256'h70352f4452351909625530004a4457331027bdbb911f0ca8f0999c9a8ea208d8"
// synthesis attribute INIT_2A of bigblock8 is "256'hdfffceb8508a8d25f3f7ff67ea95cfdfda7485e171450bce397f6b329f84626e"
// synthesis attribute INIT_2B of bigblock8 is "256'h41e7ac7a3438e4dd7201f9885a21cd606104c0297f05ffd5ffffffffffffffff"
// synthesis attribute INIT_2C of bigblock8 is "256'he9a5d488e01abb8fa350ed91729fcd366391aed58c9551a2752905b20000e440"
// synthesis attribute INIT_2D of bigblock8 is "256'haf93c73636312263115ea65c10486b4f8224fa4a719bd58b911c09f0c48d018d"
// synthesis attribute INIT_2E of bigblock8 is "256'h7274fffb9679d7ea56885cdd132dcfacef657d58ba5e31e8b22748d023893883"
// synthesis attribute INIT_2F of bigblock8 is "256'h18a14896076be067a46f5a67ad07504d2589cad219611e9899e649d603acff80"
// synthesis attribute INIT_30 of bigblock8 is "256'h1a88831be5e7f66c2526eae402fe40006c7af1e5e871e218bbeb66f49f46395d"
// synthesis attribute INIT_31 of bigblock8 is "256'hafe834e7119ad826ebaebf1e1559e2b10075d20034aab8347a59191f3cca8b30"
// synthesis attribute INIT_32 of bigblock8 is "256'h18be897109a850f365d23f87607e95fd5f2bb89eac3b88b2864fd273e366aa8e"
// synthesis attribute INIT_33 of bigblock8 is "256'hc53e92ac96b29c72ebcf26fb54bd3ac87158ebfcbf6c24586593b8f16870fab1"
// synthesis attribute INIT_34 of bigblock8 is "256'h4a3b576d1d48f2bafa1e9ae3c549af31ece5c9dbada275bf325bbf4d7ad5fb4a"
// synthesis attribute INIT_35 of bigblock8 is "256'hf464ea1ab03cc6ba58dd58b8884aae9d7feafde3ae3f5bd7e9eff623de3b07d7"
// synthesis attribute INIT_36 of bigblock8 is "256'h25378e4d09969035c62d28c914680038000062600a457199c6f3838ef37e01d8"
// synthesis attribute INIT_37 of bigblock8 is "256'h34322e06b3897d92d96c4e737c5c677a9c501e5f4a16a372a58e59614f171922"
// synthesis attribute INIT_38 of bigblock8 is "256'h415603abff807274fffb94b9967361842f43dbb714db594acc2ff086fa207b27"
// synthesis attribute INIT_39 of bigblock8 is "256'h4ee362c0210b2418641607ebe073a44f5a67595b304d1969dad2192113ea99e9"
// synthesis attribute INIT_3A of bigblock8 is "256'h03b46e1209a8623c1e5a1ddb2b3c00ede070a4200e63c8c0edb199828ddebe75"
// synthesis attribute INIT_3B of bigblock8 is "256'hffdff9dedfb78e0584478e71d94e5b08de74df347debcbadb77a83309405f34f"
// synthesis attribute INIT_3C of bigblock8 is "256'hffdff9d7be7fd35a5ffcf9ff39cf56ff0ef389768fa7db7135493fd73ebea671"
// synthesis attribute INIT_3D of bigblock8 is "256'hc8e33d3bca319eedd0daa623d3902f123e6e0a61d3a7ffff0aaaae9c89793fbc"
// synthesis attribute INIT_3E of bigblock8 is "256'h915f570e7169a5a3cafb98a539ae8e9e8021c09ac6012c2d5f14095e11e518f6"
// synthesis attribute INIT_3F of bigblock8 is "256'h44dafb057d938f8381c02347f2ae6c5b48500000d51062703695cc12ab83bc5e"
// synthesis attribute INIT_00 of bigblock9 is "256'h97ddeeded68d73f7c562223d481417ad589c281ac401d52acf59597949026bb9"
// synthesis attribute INIT_01 of bigblock9 is "256'h5ca5571ae2127ad1b874d4305db1fbb21565b513648cf29fbd596940e798771e"
// synthesis attribute INIT_02 of bigblock9 is "256'h1ec1800a15613e55040eff807274fffb2e5bd2cbf6024fcf91e786863840036c"
// synthesis attribute INIT_03 of bigblock9 is "256'hc3f446d1470f4f586d5acce4f0008b1e0f2a091587805459898d0056a63cdaa2"
// synthesis attribute INIT_04 of bigblock9 is "256'h9bf32382d3113d9ef6ebee6215b6be69b5faa41f55d755dfc3b1e0ac35a57eb3"
// synthesis attribute INIT_05 of bigblock9 is "256'h5750406604c7190fffae55ff8815d85b1e152d29998d5a99aced8b9076ac32b9"
// synthesis attribute INIT_06 of bigblock9 is "256'h7ab60cd86d099fbe1895128a30ff7d916ab2056466270a1f362a543a302a788c"
// synthesis attribute INIT_07 of bigblock9 is "256'h953d392d0c7aeb0e8935661d03e513af0d407439618f201192c661d1fc57d6ca"
// synthesis attribute INIT_08 of bigblock9 is "256'h2d6dbc5769ffca65158a03156be2a3363d3955c114b48c0eabd7fd0d36235c8c"
// synthesis attribute INIT_09 of bigblock9 is "256'h73ef38d6dedfbd9e8c413d7349f1f17e1158aded3f76d36e6b6f3cb06df68d99"
// synthesis attribute INIT_0A of bigblock9 is "256'hb4ffcd7cde3f1e9ad7ffef5abfff19cfd79799f8bb6677f1fffd6f22ba6b4ff5"
// synthesis attribute INIT_0B of bigblock9 is "256'h9deb1b17239e4a2110523ca9b8ac45241555d5ccd12801ba533b5e35ff1f5f76"
// synthesis attribute INIT_0C of bigblock9 is "256'h0010c4a4cb0235c3800216616358051dbd807074fffb276a4e342d15102a6039"
// synthesis attribute INIT_0D of bigblock9 is "256'h00281840d351252cc994412acbfd803427a690000b928b6c08988780603db157"
// synthesis attribute INIT_0E of bigblock9 is "256'h1b8c656e7f1314dffc8e0b375ba468da2e6c0e67b50829f9aec9432d7bae0396"
// synthesis attribute INIT_0F of bigblock9 is "256'h51b7e623f75e28265fde704ae8cfa1c6c8017c44243132204687e16ebef8113a"
// synthesis attribute INIT_10 of bigblock9 is "256'h0c2c0194347f644f4309949ba7eb47620bff383f12e323d9eedb8d7aeed2e28d"
// synthesis attribute INIT_11 of bigblock9 is "256'h9802544c0222822f45233955998bb33f488ad63c547cfade1086ccf68db4a8e3"
// synthesis attribute INIT_12 of bigblock9 is "256'h69adff845e11ef76ea62bc51a91c4229090113aa688e71b8cb8fcb4b78eb4dde"
// synthesis attribute INIT_13 of bigblock9 is "256'h64fcdd6ce31ffcfa23b3a78a953782eaeb3d0913bd078d9f1d23bf92ca0e4989"
// synthesis attribute INIT_14 of bigblock9 is "256'h426e128c98109d7c5bb5f9c2a8cb7ff50331e7eddd68fe7e939fa92a1ffea7f0"
// synthesis attribute INIT_15 of bigblock9 is "256'ha12386da07d2000b6080470c2ecd6f737f5cad6e7ec483e3b637729d4f6e48db"
// synthesis attribute INIT_16 of bigblock9 is "256'h70c8a61835770c3d251abd0102db8a1e232e5de9204b80037485fb726bff1141"
// synthesis attribute INIT_17 of bigblock9 is "256'h9ee3c25c98f89a7de4d5084100ce7f3be244e1880a3558c468f0030c6ee8648b"
// synthesis attribute INIT_18 of bigblock9 is "256'hd6cac95d1790670792ba228531de7cb2921716a651a60bb674f422b7ae62cc3a"
// synthesis attribute INIT_19 of bigblock9 is "256'h6e471889d5f4f6249171642a9d964eaba6fb767b9c8ba4998fd75d8c45f5df51"
// synthesis attribute INIT_1A of bigblock9 is "256'hd72531a5cb0806b20010a10d380a034f8896fbab7255bb45751be84504121bbe"
// synthesis attribute INIT_1B of bigblock9 is "256'hcf4cf72971378c1b10d0a0449adc289afeb8da7f362ce44ecbab926123845dcd"
// synthesis attribute INIT_1C of bigblock9 is "256'hfccb767f932966bbdab90720185450e39b9041f4a10cb3ee1ab969e9fc1b7395"
// synthesis attribute INIT_1D of bigblock9 is "256'h10c9a5f3723782dc18226ae0479d8b0116145d1692d9ced9a659a0e501193e43"
// synthesis attribute INIT_1E of bigblock9 is "256'h2436f5b4673ce365a1a151e7004fc000db42ce8aa9742a796155214d835ddc7f"
// synthesis attribute INIT_1F of bigblock9 is "256'hfb7223ff59ad31b78e26714408aa666787436448940baae7c96152e0acbfd32f"
// synthesis attribute INIT_20 of bigblock9 is "256'h130caea8668a16e04499e1754c582302a700c23b0a16c82fdd38175b00037492"
// synthesis attribute INIT_21 of bigblock9 is "256'ha1f165a7fbfed5fc2f104fea002ef42be2cc6cee34ecb8e21f99310d4463a13b"
// synthesis attribute INIT_22 of bigblock9 is "256'hb4db9202399dc1f4aae4923780dc323fda8b174e7faad36e11fada69f4274d1b"
// synthesis attribute INIT_23 of bigblock9 is "256'h68e58f4250b068971521cba04d26584a053c0000a608c812040e9d338a0c823a"
// synthesis attribute INIT_24 of bigblock9 is "256'h590f245a544f2ba2ba9bd7cac80f314d01f78e573f1c3c603ee54f19879d1488"
// synthesis attribute INIT_25 of bigblock9 is "256'h9a80825eb19c1c74eb934161a5ffd57f05a8e9c4167b330c0b63f8d297618c77"
// synthesis attribute INIT_26 of bigblock9 is "256'h03e6d503554ce9cd99d1ce05857a650f7dc6b8e30011040093d0b2c0ec94cfd9"
// synthesis attribute INIT_27 of bigblock9 is "256'h31eb6738ea512eeb6946e4af312a2a120d484c915c0c026794405404d8d66f85"
// synthesis attribute INIT_28 of bigblock9 is "256'h5ccaad6d5c11b65b0fe072916f980a476d9d0e963840c02c8ae06d118904330b"
// synthesis attribute INIT_29 of bigblock9 is "256'hf95f000274a2fb72efff7568df0f3e15c8acc36ab7b4d3f5effe33edbec1aab2"
// synthesis attribute INIT_2A of bigblock9 is "256'hea17cff769fe130cade86c8ab6c0e498f96e0ba4030c7301a23bd018862c5bb9"
// synthesis attribute INIT_2B of bigblock9 is "256'h8635d9d028165890c786f45e2ad88f4737d25ef6643408e9371b4161004299ac"
// synthesis attribute INIT_2C of bigblock9 is "256'hce43b4853e41c1ca5192ec0c991243a21869070ee6cac0e54949cc0c68cfb1c0"
// synthesis attribute INIT_2D of bigblock9 is "256'ha4954ffa6f560904cc15a339d9ea0487423a95e9b7c4418a7c86b93671a52a57"
// synthesis attribute INIT_2E of bigblock9 is "256'h91b9a4db000480829c8b2e6124cf4f339eba3f622c142b0fcff4b7d6866a57b1"
// synthesis attribute INIT_2F of bigblock9 is "256'h58cf208c3259c5073bf64f3beeeaaa0e840a76903e845a3af953b6b174213035"
// synthesis attribute INIT_30 of bigblock9 is "256'he4cabc974c08112cc48588f8795b244863909eda8f1acb849b042d1420c88350"
// synthesis attribute INIT_31 of bigblock9 is "256'h5bf97a06a9931fdc6acc955987ddee2c8d6c5cdcfcb44ca64b329908d1eb5f2b"
// synthesis attribute INIT_32 of bigblock9 is "256'h61aadb786dd63651be681d9e0fc145446766206316aee33464feb279d057fbeb"
// synthesis attribute INIT_33 of bigblock9 is "256'h2a22c316ddd0d44d000274b5fb7070ff5a0b454e236538883772a0c59c41e4c2"
// synthesis attribute INIT_34 of bigblock9 is "256'hdd916c1b5a95dd845ca8606830886ef4a594584043140b770a79622cba04629b"
// synthesis attribute INIT_35 of bigblock9 is "256'h028932413c5e66706c1d34592ab7551f0548845212e9994c473c42ec047b12ca"
// synthesis attribute INIT_36 of bigblock9 is "256'hbb469c2cd12961a15be7a2ac4f6cd8627d858c776d65247a8b38b7166225546e"
// synthesis attribute INIT_37 of bigblock9 is "256'h6fb338dbde4d003153babe9fea1812d53665978b32c567a1320db7abf9ea0adb"
// synthesis attribute INIT_38 of bigblock9 is "256'h03eb5535baa9ec5a7995fcf70f3702155d8dda6cc11d9c03f18254645b5b5905"
// synthesis attribute INIT_39 of bigblock9 is "256'hfef148ea2c5a46944df41115798dd922dbea4a511572fa4020389692d4686c12"
// synthesis attribute INIT_3A of bigblock9 is "256'h9b55cfcb2641fc907a9d12675975fbf3e201ed15ca1bfea0cd32c78d09448092"
// synthesis attribute INIT_3B of bigblock9 is "256'hdd1552c12a74202eda9238db9b4e9fbef572f5913635d69655d6dacdfad50b13"
// synthesis attribute INIT_3C of bigblock9 is "256'h69ddb45d024426d8a0671e6176112cafaf128ebbd93e78c6940796a584b69e8a"
// synthesis attribute INIT_3D of bigblock9 is "256'h060a00621bca2a452f0868c9425e02afc2807274fffb04917712806c140f0c4b"
// synthesis attribute INIT_3E of bigblock9 is "256'h71cd41fb83561ea6b4790b58f11aab32dda99d382821136fa09f24ab794364dd"
// synthesis attribute INIT_3F of bigblock9 is "256'h000ca761beb838161d939fc847292c70bad9e55bffdafd4b2d6326f44dff872f"
// synthesis attribute INIT_00 of bigblockA is "256'h36df2b9a342537e3f866e4ce5a0c796ed866c45eff687d59a9bbd5efdea8c3af"
// synthesis attribute INIT_01 of bigblockA is "256'h59e749c1a7567f75b3ee03b066a81dda2b32aaa3f747fa945f376381d260c78d"
// synthesis attribute INIT_02 of bigblockA is "256'hcd2a16de5d6c2a6bb54d91eb16c741629f124f88da0124b4368a124ac286ead5"
// synthesis attribute INIT_03 of bigblockA is "256'hfcb280ccca51f7ff2c9c36573bb6791be6fe194800e780a3e3dc15e52624ccb7"
// synthesis attribute INIT_04 of bigblockA is "256'hc89ebabef9f339d4cab41f79f6f483ca7dd485250dfe3f512995adf68809b1d2"
// synthesis attribute INIT_05 of bigblockA is "256'h500dfaf245b208888d1fcbed18c016d46d55475b522692046fc34324796615fc"
// synthesis attribute INIT_06 of bigblockA is "256'h0a2e0003469e89232f983688cb4e5194c91a68b1d08a1ddaebd45109966f94ae"
// synthesis attribute INIT_07 of bigblockA is "256'h18b875a67907088b0105ec2a2884432868c92d5e027cd0007274fffb80a65d77"
// synthesis attribute INIT_08 of bigblockA is "256'h63a5830c0ecddba315ccb42dfb1bd516c8cb2ecd720577f221f1b461136f80b5"
// synthesis attribute INIT_09 of bigblockA is "256'h5550d022289e6f767a70fbe5c7fb3b7f6ffafff48dfebd0a03d9c23e889796d2"
// synthesis attribute INIT_0A of bigblockA is "256'h284757ed214c557e9755523532d833c4f3986bb54723519289a4ce11c1811921"
// synthesis attribute INIT_0B of bigblockA is "256'he4fe5d852f13e0696138b1d23bfe90002008c6992a42a400013eccf9ef2e5b1f"
// synthesis attribute INIT_0C of bigblockA is "256'habfb850b0a5ba1712c8a31c3ba4ab86829077fa33b5f64bd6aa2fad7af65fa2a"
// synthesis attribute INIT_0D of bigblockA is "256'hc51671d7aa872080a0d6ec8bfa3e23e9ffb3d3d1e31fa9bfedfa18347a7bddc3"
// synthesis attribute INIT_0E of bigblockA is "256'h51d99ccb2255ae86a559214f08db94a10ccd4f88887746d7226eb6881f87c959"
// synthesis attribute INIT_0F of bigblockA is "256'h4336241d8442213cc8101c554890e30265a8e1f880ec06feaca696c030992c4f"
// synthesis attribute INIT_10 of bigblockA is "256'hfffb47570827d3c2e3c12b8822da71d7399bf9706d9b272583ecb0b61031186d"
// synthesis attribute INIT_11 of bigblockA is "256'hb41390ef209824567da335330c4a0062dbed280415ba6926585e0312da807274"
// synthesis attribute INIT_12 of bigblockA is "256'h0495e6aa4e8e7d3f7f64ed3307efbf7dfeb11811aa8d4eed8be04b78c2600858"
// synthesis attribute INIT_13 of bigblockA is "256'h5bf40d3454428374b683eedf0bb80b12686edafc2ec60248d400f5002d9dd03f"
// synthesis attribute INIT_14 of bigblockA is "256'hc5388980a1a0e50f488117040220cb3319e5dd4cdc901adfdb0aa5a2f5f9dea5"
// synthesis attribute INIT_15 of bigblockA is "256'h341232feb9a5d4f1559998e368e72d9e2bb1fdb47b63fc4fe0843c90824d8951"
// synthesis attribute INIT_16 of bigblockA is "256'h46bf29b70c315f33879e475f1aee23ead58dfa02a434cc0296ad47e6d630efe3"
// synthesis attribute INIT_17 of bigblockA is "256'ha03db100291791d5bb2d566ae39f0a0d89e5b565118d8022cf5c3f663a755b46"
// synthesis attribute INIT_18 of bigblockA is "256'h178dc29640e2a0468848407320955d81dd8116fbf121d43af52c10f4884a4f72"
// synthesis attribute INIT_19 of bigblockA is "256'ha9e31876ec4956b3e7dcd42dc04753b89d5bcf4c999a80b75427dcc7a1388cd8"
// synthesis attribute INIT_1A of bigblockA is "256'h02c1e4807074fffb0da59e169a313d5d8c183db7301c41de74f9f1f0b789e225"
// synthesis attribute INIT_1B of bigblockA is "256'h89fa1fa119b8b481946ee0af945875445535080a01221baa2b652bc8698b4d5d"
// synthesis attribute INIT_1C of bigblockA is "256'hb69f2512ea1a99951ea1f56be10bffff12ec00009ff5e06f22ca5ddb48223052"
// synthesis attribute INIT_1D of bigblockA is "256'h05e6dde3000644801282683fefcbe221b6e5f5104d466aedbb44f6edf614b436"
// synthesis attribute INIT_1E of bigblockA is "256'h93f6850091e9d68b491fb5469efa467253a766e37aa3a584e8a1431ba477d150"
// synthesis attribute INIT_1F of bigblockA is "256'h2fd9ac47a4e6ae794169fe712a236b38e6ed5d83ba90086f7dbd9bb975ea98fd"
// synthesis attribute INIT_20 of bigblockA is "256'he917ffa20817ff20ffffffffffffbffffe9a05907774e5f7dcb665dada3f3d3f"
// synthesis attribute INIT_21 of bigblockA is "256'hd401186a8554dd1db7b8ff2f465e263dc8f3af4124d85a619c511a4ea31b0348"
// synthesis attribute INIT_22 of bigblockA is "256'haa5d36659e127ab05dc6e2eb46796c36c8ddce0796706f0bb13111cfab1344cb"
// synthesis attribute INIT_23 of bigblockA is "256'hf0e27f58848795045e622f43906030d2cad7728609bad48aefc9c62c1764dae2"
// synthesis attribute INIT_24 of bigblockA is "256'h3829272e5bb1b64d000274eefb72fbff6f722c6ffcf61f55554f674909d3ba23"
// synthesis attribute INIT_25 of bigblockA is "256'h8d77009b004053e88e7e38b293156de4ab94ba60c49c096e4ad1050e7701e4db"
// synthesis attribute INIT_26 of bigblockA is "256'h71d02f2330fd53a7d3e7f91f657a7432219b5961ef0747be4fb90c76f0f472f2"
// synthesis attribute INIT_27 of bigblockA is "256'h2bd5d818eb6506809cb4579670c2a69c11fd588e346c2d1f019c19500200c3b2"
// synthesis attribute INIT_28 of bigblockA is "256'hdf7677c7ac28a57364ceaba2d41feb530e73f4e10eff44c63768773e581e7ebd"
// synthesis attribute INIT_29 of bigblockA is "256'h5ffebe8f39da7548c1b12d6b30b753f6dc216d9e7602170990d2ec5026d42c1b"
// synthesis attribute INIT_2A of bigblockA is "256'h6e47282d7711d9d0f9038b18a8cded0bfcf6fff04a8938b12ea51ae401490801"
// synthesis attribute INIT_2B of bigblockA is "256'h70a381f3384f45492a4ecb9783630a4802ca400172a04c876f17e5e7b7b6dcb5"
// synthesis attribute INIT_2C of bigblockA is "256'h9e6b689b45722d1a90beeebcfc8689a61b7cb9acf7d46152b9dd942b369b8a90"
// synthesis attribute INIT_2D of bigblockA is "256'h29bfa9e528ff971f9c6d109b9994e39c5b62a4f1c83f2009f368bf42890b3587"
// synthesis attribute INIT_2E of bigblockA is "256'hc20e660044dbb8258b54db391047000374f8fb72ccff6cafd27ba617ac3ea8c5"
// synthesis attribute INIT_2F of bigblockA is "256'h8d6748d2034c19d1c63d36d70a0a04001980619e6d9ca013fa60a6141f6c0af9"
// synthesis attribute INIT_30 of bigblockA is "256'h00130402062933947fb8bd4d9e7e9dfab323da837261289e47ba9e1e7e210a67"
// synthesis attribute INIT_31 of bigblockA is "256'h96231af9f5223f9798cae24861a8a213359ef6c570ac7c7e17ba519581ad75c5"
// synthesis attribute INIT_32 of bigblockA is "256'h5453f59874e64060b3cd3f514171b69d792dcd5efa3513a027163199fc274358"
// synthesis attribute INIT_33 of bigblockA is "256'h28e34020ffc0d5ff6ebb3147876717959fe89a0218bf6ac28365007661769c41"
// synthesis attribute INIT_34 of bigblockA is "256'h8e90feaf3bd9009f00bc64c528dbb48b35554f8b9a1d8c2b01c84a2710d35db6"
// synthesis attribute INIT_35 of bigblockA is "256'h243d790f624ae4c73ae43aa363e364a319aac905a4ae0400a801c1dc9dc4995c"
// synthesis attribute INIT_36 of bigblockA is "256'he27f219a8d64809eeebc0593b38a00c6bc08906d28c6e7ebf58a8647aadd6d2a"
// synthesis attribute INIT_37 of bigblockA is "256'h1c4fad669bc98c7dfa0fa59b59fac48bea881e50b1fa709cfe446e2f50603197"
// synthesis attribute INIT_38 of bigblockA is "256'hc4a01d6a0bf9270e5701851ba82b8716dac9ef46800274fffb7200ff53fd15d1"
// synthesis attribute INIT_39 of bigblockA is "256'ha5d121c572b9ef79d54f992fe8dc890431825dd3a36d609262a26d68b393f8a0"
// synthesis attribute INIT_3A of bigblockA is "256'h0bc9279cb45a0cb00490103050af292837aef8612ee8dbb3b584a703aca2c326"
// synthesis attribute INIT_3B of bigblockA is "256'h70e7053fb7bd35beeed15c12869d4c6e6a5fe168ad7cb41465fb6de56a09e281"
// synthesis attribute INIT_3C of bigblockA is "256'hbfa477fd9cc31f2669ffe503ce2d83e7938a6ad27ca5657c8d33f8e00d1ce837"
// synthesis attribute INIT_3D of bigblockA is "256'h216a559e830b248ed669425c5b47577e71b82004e020ffffffffecf4efaf1bbc"
// synthesis attribute INIT_3E of bigblockA is "256'h4a6405222001dbd2df408cd747cac7a7f1fd0c4d8e267920b67fd72a6fb8a292"
// synthesis attribute INIT_3F of bigblockA is "256'h00b59be67426162293d6c26f5d4549b4c2f8a2a5bc366c5cda15bcfc85d7e594"
// synthesis attribute INIT_00 of bigblockB is "256'h48c8cf6326bac5625d513752da1c9ea7226d3e40e7a92191c4d6391d5be48009"
// synthesis attribute INIT_01 of bigblockB is "256'h00ff800825bec8abcb12444df7cd7457c24bde71a9975931663a301427361a5d"
// synthesis attribute INIT_02 of bigblockB is "256'h6d4cb2945660c6191d6a0bb967785718651b382b8a16dab1fa47800274fffb70"
// synthesis attribute INIT_03 of bigblockB is "256'h50193753e14b36956759050710cf1404921d02af5c6559741af700b728099116"
// synthesis attribute INIT_04 of bigblockB is "256'h7314cff593eeb2328a702486a167a78d95578a10622a124ac9d0b3b64b74904b"
// synthesis attribute INIT_05 of bigblockB is "256'h048eed82d4e582a8d027dc7c13a8ef9774175a8522e1ec79cee13f2c9b381330"
// synthesis attribute INIT_06 of bigblockB is "256'h7fa6852bfce2cbfce7df6a32c2fb4c6da5af9d0a1bddf881a35700f4ddeb0c79"
// synthesis attribute INIT_07 of bigblockB is "256'hff86e2efdd378e93f8f49b5e6b3affebe3760c6bda625f5bcdab297bfc5d358c"
// synthesis attribute INIT_08 of bigblockB is "256'h50d8b19e2606252c5c6a18b26443ed1dae4046dac00099f4a6bffd76e7efa8ff"
// synthesis attribute INIT_09 of bigblockB is "256'hd5bccffa93fd7ce9656d4d09c4a08ad79bdfeec1a97b2b901f919b6a04ce0cef"
// synthesis attribute INIT_0A of bigblockB is "256'h04a91157e49758bbf578d0b130b968c4d4ad75279c8c4e8891e500000000535f"
// synthesis attribute INIT_0B of bigblockB is "256'h02abff807274fffb2b0a95d32b221711c689759eb1588ea3c54e8290da5a10f1"
// synthesis attribute INIT_0C of bigblockB is "256'h8b4b1cb615682894136d20ba255168465537c00c2447db472f841630318741da"
// synthesis attribute INIT_0D of bigblockB is "256'h2e5c84315d92d572d0f79521d8356f8f144d30dc0d51cefe895fa6a67c6591c7"
// synthesis attribute INIT_0E of bigblockB is "256'hfdadf4791af77de76d668ac1816c2469110eb8231dcfeedb67c7edd355b810c2"
// synthesis attribute INIT_0F of bigblockB is "256'h1fffe0e00b83e800fd16bae583ae18ba07f0fffeffbf7f07727fb0647162cb82"
// synthesis attribute INIT_10 of bigblockB is "256'h5299d133c735948d1c1851fa2ac525d74cace54085225dd0c2ded12ec24bffff"
// synthesis attribute INIT_11 of bigblockB is "256'h59ca5bb8a8745b2db496ca6e91560913f33de4e0e96c22d1f12432c397c769b3"
// synthesis attribute INIT_12 of bigblockB is "256'h1f0e19ad1ca82c3ec25c0e9bf8623ec1d990783db72d95c0a854bcfa84ec7242"
// synthesis attribute INIT_13 of bigblockB is "256'h1edcea963d5e253a2e5e67b2172f72ac36d19e9cf2cadea19350075279069f40"
// synthesis attribute INIT_14 of bigblockB is "256'hb5acf6e5448e8eb54abe2a27b454e78cc95fc7482a14b321ada276b0403bf04e"
// synthesis attribute INIT_15 of bigblockB is "256'he008853d4cd803daff807274fffb3fecba6fbd2b516e71fab547f50d72965aed"
// synthesis attribute INIT_16 of bigblockB is "256'h7bf9d7ac9bb95e66396ac0004b1e8f2c00f587806259ed190052a624db133804"
// synthesis attribute INIT_17 of bigblockB is "256'hffff0080ff00dfcea266497f666b7d2663ebf46a66fdffa68d6da6d2ff36065a"
// synthesis attribute INIT_18 of bigblockB is "256'hd68d1a9c6e6c7695d87d445648d17998309117402f2dd324330662237260fffe"
// synthesis attribute INIT_19 of bigblockB is "256'h9fd565bdab446915a714cf544bc0000d204014d0129c228e455f55d7f5b44156"
// synthesis attribute INIT_1A of bigblockB is "256'h9dab0b60cb554b31189c800b5912bd9d92aef7c689c7ed909eb03221cf509603"
// synthesis attribute INIT_1B of bigblockB is "256'h1da19d2c0fd261741b0146fcc4b5d99a45e0e2574757af374ba8b197bd47fadb"
// synthesis attribute INIT_1C of bigblockB is "256'h1e8ee77a5fe874bd3fa7b177e6f73aa4ee528fec8da3639012204fd66df7149a"
// synthesis attribute INIT_1D of bigblockB is "256'h1fffc0804c636633b3b1e4de5dbaa6e6d4ed7a69fe98dd7cede6696bf48ef93d"
// synthesis attribute INIT_1E of bigblockB is "256'ha582109d56fdb1e67ef805ab7e6afd3fbd5b909459a221d843a15255d933cf07"
// synthesis attribute INIT_1F of bigblockB is "256'hc624cb46328380000661645a04e0c6807274fffb0864ec42e41e2935b8485475"
// synthesis attribute INIT_20 of bigblockB is "256'h6447ef55f72459619419cd6446b0e86e90011b900b6d208bf60068dcd9830011"
// synthesis attribute INIT_21 of bigblockB is "256'h1cbd47b97db5a32e91f5a9003779144b2a9c69b1b4bba0f7f4e0355c8e612372"
// synthesis attribute INIT_22 of bigblockB is "256'h40bcdeba57ab2b27ddfff79d3bd9066e15d069cea73f80145b25573bdafe8fa8"
// synthesis attribute INIT_23 of bigblockB is "256'h991a22446016d50cdc6bb33ab6170c4c7f0975345faadb44d8e1f74cb4d6e46d"
// synthesis attribute INIT_24 of bigblockB is "256'hbf1c981c07a39fd3f9900c8f368a0c1f30b9156c3a46a55348126a4245406536"
// synthesis attribute INIT_25 of bigblockB is "256'hcaeb59aaae6556a951ee59244a54ea9e9a03de314adf9a20959a0248503d8b3d"
// synthesis attribute INIT_26 of bigblockB is "256'h0439e8610969d1102a26a2a24a48342736360a0b439b3abc6865bbe5f79432cb"
// synthesis attribute INIT_27 of bigblockB is "256'h2652ab706fad9e0ce0518e8fccf373d059cf1e09b3871480c7dd209b255f236d"
// synthesis attribute INIT_28 of bigblockB is "256'hb87f521dddcb722586afd32f044d562468fb09bbab95a28860ca4ad5532e2d4f"
// synthesis attribute INIT_29 of bigblockB is "256'h75a34d072c4c04651ba71b831622512341dd02dc91807074fffbebdaca2d5b0e"
// synthesis attribute INIT_2A of bigblockB is "256'he6e6a596efbf727a48ad6581d0c8821d9b5eb2799fec99d0a8518dee40822055"
// synthesis attribute INIT_2B of bigblockB is "256'h28640e1557657e930c28d5bf5dfc91374a9f0be3fda33212f5b34368faea3a99"
// synthesis attribute INIT_2C of bigblockB is "256'hbfb5acbed40fd7125bd7925e902342db8b705cef63b704e94909c8db062f6288"
// synthesis attribute INIT_2D of bigblockB is "256'h46d793f345868719cc28090fd8bda98e3da74e28889ceba7a180451236b42c50"
// synthesis attribute INIT_2E of bigblockB is "256'h49874f9308c8bbf7abf0480eeafff556f7ab6e6afe8502591dc9a80f00859239"
// synthesis attribute INIT_2F of bigblockB is "256'h734a0d87d53bc546d3c2a235449fa262b93ae95c6843ffb924f552e776de56d6"
// synthesis attribute INIT_30 of bigblockB is "256'h10c42beb2cfa299caabc70078f9cb3621afd9148161617832b9a1b6d7b5934c2"
// synthesis attribute INIT_31 of bigblockB is "256'ha0f89acfa475644c3a0b33f0bc956939c156a8cd8c6aa15218a8002024820401"
// synthesis attribute INIT_32 of bigblockB is "256'hb9ff31ee761e9f4068b9846de4cf4f3fb71195e6ea28f2b7e1560550d58cae1e"
// synthesis attribute INIT_33 of bigblockB is "256'hefb4830d6fe0a6200b790bf12874ef18e2db2220cc2dde68e7470002749ffb72"
// synthesis attribute INIT_34 of bigblockB is "256'h53debca4d727f2bc4a69452b94569a1c25be6fde6bcdcbd7710a97d808823095"
// synthesis attribute INIT_35 of bigblockB is "256'hee316f0c72b4509194363af7554c8ce56d04c923000d018049e12d09d0e24769"
// synthesis attribute INIT_36 of bigblockB is "256'h71b713d67b0a3e9edd19b0ef585c4c1a59611e10c1b7890b42921b2001994400"
// synthesis attribute INIT_37 of bigblockB is "256'he3ea0fea1351256aa41404fae691ae58a3e777d17e9c92aa93ebbe50ce23605e"
// synthesis attribute INIT_38 of bigblockB is "256'h0200086bb1615448709cb51eafd463a141e1c6847eb2d0e3236f4dfe9a366444"
// synthesis attribute INIT_39 of bigblockB is "256'h100004006b08f983af044fbc0b1a955f71a70ad79f5189953583a7638db414d3"
// synthesis attribute INIT_3A of bigblockB is "256'h9bff5dfbc6423f9d294a4c45a3845939422a3686d0385dc8688c8e502da425d8"
// synthesis attribute INIT_3B of bigblockB is "256'hb57f74ca22f57f90345d1b7ed87fbf54006ab180be835c7241dd2b11a8482447"
// synthesis attribute INIT_3C of bigblockB is "256'h000374abfb7200ff56420045ebc467b4d16965249d079b55dd15e9faf5abfabf"
// synthesis attribute INIT_3D of bigblockB is "256'h05724800238a6e28750cb6e044a00b710c1d63068d0ca1cb2a15272edc69225d"
// synthesis attribute INIT_3E of bigblockB is "256'h3735cfac8c6efda7b5601d850000491981c607becb9435648424c830495136dc"
// synthesis attribute INIT_3F of bigblockB is "256'h716ace83608c2ca28608568aed68475b904be39014671fce02ce44b3e0e4bc2b"
// synthesis attribute INIT_00 of bigblockC is "256'h70e9479fc5da5c54b5b6f9e2d1cd94407cae6660cc0fd4b2c9b680802389bcf4"
// synthesis attribute INIT_01 of bigblockC is "256'h00008800ee1ec1e792edffa2ef3fe62f0879c3651ec559ce6bed7ddaffc5ff93"
// synthesis attribute INIT_02 of bigblockC is "256'h96a352243d64436549b620899188e5a9bed1f9a351aa32060c83459c2369b249"
// synthesis attribute INIT_03 of bigblockC is "256'hbe154e3a7e759a4cd82ffab7c1b7f56370d7932e41c962c339f14598ae3e5dd7"
// synthesis attribute INIT_04 of bigblockC is "256'h54bad49fe7ff28fb6459918562dda86c63d8507e0eb34bd0d9d517ab3f84a8fe"
// synthesis attribute INIT_05 of bigblockC is "256'hc88146daa59220a0b10802104c94a40928b95fcc4acb49707b76cab4bd2821e4"
// synthesis attribute INIT_06 of bigblockC is "256'h2c2b5ad1df4f000274bafb72c1ff600deeb73105a7f8d7a0628e39306d9b2a54"
// synthesis attribute INIT_07 of bigblockC is "256'h49cca6105229a4a0904a63986d745b0678e8c61d0d6a4d6d23505d20017b5016"
// synthesis attribute INIT_08 of bigblockC is "256'h286bd49ecb943efc9538c79362589136995cb58b5d02bc0f7aaa4716c1ba84ed"
// synthesis attribute INIT_09 of bigblockC is "256'h9b65fd29badfe4b4244d4ca065f850cd9ecfc2d9b39406f7350a7ad1c68f1037"
// synthesis attribute INIT_0A of bigblockC is "256'h3e716da546a39c1d1ec7cfda98e4a101cd55994008c23997ba50353dc9bff0f4"
// synthesis attribute INIT_0B of bigblockC is "256'h911233881b284e644249e4012285c2f0c86404876f624a04c65b989fa0c94327"
// synthesis attribute INIT_0C of bigblockC is "256'hb1b1a1e37a5ee837a3c469001327a46e67e8b4c5631406ef2ff2414c2160931e"
// synthesis attribute INIT_0D of bigblockC is "256'h990ad80c290ea72753f45cae182f7e628dad14f5aae23ca267bfa00e302ec752"
// synthesis attribute INIT_0E of bigblockC is "256'hdb558d24808a0188daf2549a02d640be06f695d66ebeefd80830fabf658e9727"
// synthesis attribute INIT_0F of bigblockC is "256'h85902539800125801a1b4936c33381373eb5d082d0ebfc36286d484691485b1c"
// synthesis attribute INIT_10 of bigblockC is "256'had0ce2db281d2b3edd69194d000374cbfb708bffd471a996902a688eafac12b6"
// synthesis attribute INIT_11 of bigblockC is "256'h003b363467466b2ecb8b0de44cb1c0ce308c6ea8700b78a0a49433750be1463c"
// synthesis attribute INIT_12 of bigblockC is "256'h59f9e5d4eb13be82e5cc7ad685b9a3a985fbb265b7dc16ff9c7302298547062d"
// synthesis attribute INIT_13 of bigblockC is "256'hf0080ce0f4b854cf7efdcf0ec2b21d929f0193f0cf4ea7be710bfa58214bd91d"
// synthesis attribute INIT_14 of bigblockC is "256'hfdf6bcd0a8442e740b20002600208124fae169099a97f68776a4df36a77f4400"
// synthesis attribute INIT_15 of bigblockC is "256'h95ef160466cababdcbb2b70a87739fb467af23abe84be2cc90d6799b745a9132"
// synthesis attribute INIT_16 of bigblockC is "256'h9a9a0cad65ec23c572fd8b66d59134128430a9bb2899b47666d6cb8a83a72d13"
// synthesis attribute INIT_17 of bigblockC is "256'h001086ab1872f901d0b0dad32ce803940303c80366428a083c502822562399a0"
// synthesis attribute INIT_18 of bigblockC is "256'h3606a21123c581aa00010000a98134ff72953b8066d2b686ea2dd5057fff0002"
// synthesis attribute INIT_19 of bigblockC is "256'hd30cd0863480e0e7cbd4026bc43ae45eda18699255ad11cec96e2b54c7a19caa"
// synthesis attribute INIT_1A of bigblockC is "256'h71475933580c2066db8d20421eba51224ddc0324d7807274fffba68db391270e"
// synthesis attribute INIT_1B of bigblockC is "256'h6423233bff241985d98308b7769cac88c9e75101dc418d49306005eee84ea467"
// synthesis attribute INIT_1C of bigblockC is "256'h2c00c899c423581fda6ddeffd3f94fcfffe7def9579dad8ef72ce9a799a1999a"
// synthesis attribute INIT_1D of bigblockC is "256'h30764ea02c06012a0000081a828f8992782c167b7a12987d695cb49304510000"
// synthesis attribute INIT_1E of bigblockC is "256'hb0830c38a6b12114a89038b4e4080d52c2cbe60e48ba1c2cfafa4b8381737ec1"
// synthesis attribute INIT_1F of bigblockC is "256'h40afc51669c766a49fd2943934e7050ebe9d07f55b8f58a05105dc85355b51dc"
// synthesis attribute INIT_20 of bigblockC is "256'h4000a0f5daab1fcaef16f133427549abc50485bee9197bf3169166c2a666bc3f"
// synthesis attribute INIT_21 of bigblockC is "256'hc9eaa866a14cab41000ab800514b67d91b25bc42c358a46814c9dc4a97ff0000"
// synthesis attribute INIT_22 of bigblockC is "256'hbe84a32957259347d182ae2037597dd53ae1bd531c5a11954244046e41a3c372"
// synthesis attribute INIT_23 of bigblockC is "256'hcf62a39c383b9fe06ddc46b7c273a7285968b9b4fd7aa8b24e75bd43cfb8c9db"
// synthesis attribute INIT_24 of bigblockC is "256'h852d285818736ae6f565140c0526ab5c15411e18b18643da0360e5007274fffb"
// synthesis attribute INIT_25 of bigblockC is "256'h5fca4c26ee7ea7f2588238544c8bd3e229bf3b2c327638b520bc25d220517413"
// synthesis attribute INIT_26 of bigblockC is "256'h3d706172da4b2a6c707213b628a3b68f1c910037cc00a3f233b6c6174dffd4b8"
// synthesis attribute INIT_27 of bigblockC is "256'hc800d6e54b49862eaecaac0ee35228543c4c0830b9096d8f05d4920000181b02"
// synthesis attribute INIT_28 of bigblockC is "256'hdab5b6f6004735812bfbdb4a674c78b6cc7c31e609665a7b70087d41b651dae8"
// synthesis attribute INIT_29 of bigblockC is "256'h1dc9b132f9f2417e72708cf2615959fe84a47ff961ebf48a2bcf43bdc53f04eb"
// synthesis attribute INIT_2A of bigblockC is "256'h2a93a287487a19a8143667e8a069e46d049434e00fc3056ca5016513080ac251"
// synthesis attribute INIT_2B of bigblockC is "256'h1e1bbc253e504d12a924428c1730003a0102a2a05262f39090c67450167d6e41"
// synthesis attribute INIT_2C of bigblockC is "256'h387cde81f8a76d2185bf6b6c1be68c6073e7f610fb4bd633e6d149d9bb7f9cc0"
// synthesis attribute INIT_2D of bigblockC is "256'hf0807274fffb4c2116fd88e3fd9c1611dd4e97a599949988cf632f0dea78759a"
// synthesis attribute INIT_2E of bigblockC is "256'h69f69819681405ad2859147e6a664513000e0426ab5c16611d2ab9864d5a034a"
// synthesis attribute INIT_2F of bigblockC is "256'h40b407754dbe31ca74aad9b3db4525c81000d4205faf303fabeb4b047522b59c"
// synthesis attribute INIT_30 of bigblockC is "256'h4a814b64352cd2b268f14361a85d62550101c00041abb50b08656a808febb368"
// synthesis attribute INIT_31 of bigblockC is "256'h86fdf3924ea35dd1552ebbde9cf13e9bfe70ff89f6d86b6d5933a6bcda8822d2"
// synthesis attribute INIT_32 of bigblockC is "256'hc750833da2509fbaf7136ae5dc1cbb36510e188269c65aaccc0e540c99cb84b5"
// synthesis attribute INIT_33 of bigblockC is "256'hc100fffffffffffffd5f4f6fa8351bf7cc8c51a9aee16abe1214ebe73ac9da34"
// synthesis attribute INIT_34 of bigblockC is "256'hc15205eda060217d9698d9644187806b194e502cc0d300c8e5bdd685db7b2648"
// synthesis attribute INIT_35 of bigblockC is "256'h98bf7631c4a6e67a8cbcc30a49b5d459024a222bc13ea179338000450028df70"
// synthesis attribute INIT_36 of bigblockC is "256'h89413dca31f6054c2ce7be33d420397bb432aa2d1a6014e68f67238d421e5b7d"
// synthesis attribute INIT_37 of bigblockC is "256'h51264ddc0363f7807074fffb96d7e3c6e95bb77952268485d9959dadd0dba774"
// synthesis attribute INIT_38 of bigblockC is "256'hfa1bad24d42cd647083028138d6e607c99517124910d164b04c5bb871f021f18"
// synthesis attribute INIT_39 of bigblockC is "256'hcdae04c5d73e3ec99d90709af2ad7c93cf5463328747ab1888e56eadc923e800"
// synthesis attribute INIT_3A of bigblockC is "256'h79e5d1bc57c748c3568db814c7247cd96864ba509a6b6db11881100406c11f47"
// synthesis attribute INIT_3B of bigblockC is "256'h26864735d8b7d9d1977f4a4bcde296be3fa46e0bef1e5936e14a12561deccff2"
// synthesis attribute INIT_3C of bigblockC is "256'h4a0ebee23eac7dfcce19df1bab3fe6f6c6dbebb17b6d734d68efc973c87da19e"
// synthesis attribute INIT_3D of bigblockC is "256'h9a67625965c7a4d4dbac724800c1fffefffffffffffffffffffff57fd1e974a7"
// synthesis attribute INIT_3E of bigblockC is "256'hc0b23282549a003682080f40966910e14a3f1371b3c193024f4d821579fef607"
// synthesis attribute INIT_3F of bigblockC is "256'h37517214cda83616adb5c6d763ae4d5b6addaeaf48f61c7ea7850df4fcfa03f1"
// synthesis attribute INIT_00 of bigblockD is "256'h0a8e3b50df9ba21fae0cbdcd083556c1e26d091fd58ad7d9ce4a7a442c5b3adf"
// synthesis attribute INIT_01 of bigblockD is "256'h5730231b4823eb16dac1924d800374fefb72e4ffd38c2e9c38a08fa76d103488"
// synthesis attribute INIT_02 of bigblockD is "256'h6dcaa92410a0dbe9cfa3aff8ea3e5163b1966d4c8c0df140e6240f6a4b75a346"
// synthesis attribute INIT_03 of bigblockD is "256'h04400ac8c8e844ba94b12a57e569672993c85a1bd9c3cb343697322a78a86824"
// synthesis attribute INIT_04 of bigblockD is "256'hb8dce677e4245cbce9938519949512e5813f7703136200e284d9788406209000"
// synthesis attribute INIT_05 of bigblockD is "256'hb22b201bdbf0c4dd95178a237fa9f7aad9c395d4ddeb52e5d490df9b89136b82"
// synthesis attribute INIT_06 of bigblockD is "256'h03f6d44e44c9a69e4536c60f5ae371599b8e4b6a5e6f8a21e816c9b1fdcfc61e"
// synthesis attribute INIT_07 of bigblockD is "256'hf69b58f6ae11f79c5b3d8f1f18080f9961486e6429240008f810bb554ebdfe82"
// synthesis attribute INIT_08 of bigblockD is "256'hc19d8ea772173584919a0fd6898f0000002c00e00354b39985c2970c53906429"
// synthesis attribute INIT_09 of bigblockD is "256'hd3b955239713075047711dbd01a25798fe8a1eb454498b4bab04c12f0496b1d4"
// synthesis attribute INIT_0A of bigblockD is "256'h8c353d2e14a1728a506ddacff35e7bfe0a35e62eb856ac1baf806d4e3fc3fc48"
// synthesis attribute INIT_0B of bigblockD is "256'h376c4c0d46946724c35bf8238959db416f43800374fffb729affd291409ae74e"
// synthesis attribute INIT_0C of bigblockD is "256'hcecc238dc8258300df4b478b7a6de4142a1cdce0388e04946d9c900db720c62c"
// synthesis attribute INIT_0D of bigblockD is "256'h00201ff3cf7db375282e37f90991133d592a139229062ed0091921e060127485"
// synthesis attribute INIT_0E of bigblockD is "256'h9977efd64869aebddd85e3c7e0512b901937a243951129294ed368ce06eba000"
// synthesis attribute INIT_0F of bigblockD is "256'h1396f3240d5ce5d7c292a5bdcbce9b1bd678b3ab273ecae54fe395676aa66729"
// synthesis attribute INIT_10 of bigblockD is "256'hbcbb86faea86032c04de4c95d1185cb4f55ae2f3451fa0639f5bf6fbb4b1d973"
// synthesis attribute INIT_11 of bigblockD is "256'h7a05e8098e597b9a82341baef6cb383c4d6cfc9691c900a4fc104c1bc30590f8"
// synthesis attribute INIT_12 of bigblockD is "256'h76e4d10412d3b7269dc0211789d1bc38d4aa257400060010aab21ce2ba637349"
// synthesis attribute INIT_13 of bigblockD is "256'h5deec192f35dbd53322f8de57f7994cc7e96d0dd7a02bd80d61e6eb5ddf268e6"
// synthesis attribute INIT_14 of bigblockD is "256'hcda31d2a7a3204496de450e76e483955bb14b13c793528db86e67b2da38862a1"
// synthesis attribute INIT_15 of bigblockD is "256'h928db1e046240d6d0d31c2766a24433bb8252b45db394543800374fffb72daff"
// synthesis attribute INIT_16 of bigblockD is "256'hc2eee0bb296692571923900031c867929ae7146cdcdb4835e99f4985609a6d9c"
// synthesis attribute INIT_17 of bigblockD is "256'h7294903200c4120053a834550b486626c4686ee7aa60c0b1388b23913f9157e8"
// synthesis attribute INIT_18 of bigblockD is "256'hee13708170feef2bfbfe987fe3bfad1816403f7b283098559218662c2534f3f2"
// synthesis attribute INIT_19 of bigblockD is "256'ha3bb1060840a2eec40681c03e8281a7bfbf0944ddc1ce25d9f2375b9f3112499"
// synthesis attribute INIT_1A of bigblockD is "256'h6bde764fced910650408cef54dbb73c25d883bdcc5fcd53ebbbb521fbba7c705"
// synthesis attribute INIT_1B of bigblockD is "256'hdb4472463aa401447df632721bc1db994509d93a143040188324213ef6bcbb2e"
// synthesis attribute INIT_1C of bigblockD is "256'hdddeab31febb4961fad5280d005d486488d4c11251102b43fe4d293e2c72a27d"
// synthesis attribute INIT_1D of bigblockD is "256'hb93e3bbcfee99f05987794f90b41e753716ebfde26c69d5d79ddbdbd2b85530b"
// synthesis attribute INIT_1E of bigblockD is "256'h74fcfb7045ff3e4ee5b799956f0fbfd8cbb2f33b39319333ccfff48b98eeaf8f"
// synthesis attribute INIT_1F of bigblockD is "256'hd043c1892d9c840d4de0e625236c0d2122946724435bc8208b2d5b3946438003"
// synthesis attribute INIT_20 of bigblockD is "256'hbbf2268a3c5c1971b45a5dbceb9c8e8459d7303d62495e3ef7c3e5d2d64eccde"
// synthesis attribute INIT_21 of bigblockD is "256'h3130012519ba07d46076ae3718d240f91801428bd76b6db6c723aba51c169552"
// synthesis attribute INIT_22 of bigblockD is "256'h8eac0e35091a5dbb2a81760ddbb930aa51cc8638c71df7e2b5c9f78452e2dbe2"
// synthesis attribute INIT_23 of bigblockD is "256'hf7ff9145b4213b14fb5e67b13159da2457d1e287b3be37207d983c918902e81d"
// synthesis attribute INIT_24 of bigblockD is "256'h01622d5fa29876df4a3f37fddc75936e415711ead317ec650d61dabf76cffd54"
// synthesis attribute INIT_25 of bigblockD is "256'h45047190cef4258029f326463f1f2b826ab3f22da48a25e1da356da527230001"
// synthesis attribute INIT_26 of bigblockD is "256'h0477119cdda2dd20e73063a18378c6b1f3d7ad591cc0274baf8a40008235360e"
// synthesis attribute INIT_27 of bigblockD is "256'hac8ae6b625e15b1a03fe4a593ea0f16dc58fad26695f9c374e614144b1809032"
// synthesis attribute INIT_28 of bigblockD is "256'hd18860de0414fd807274fffbe84fc316f415352f1fcf3175239536319d1ffe73"
// synthesis attribute INIT_29 of bigblockD is "256'h87dc2ec28235a9b90c58741306afe055b0c17ba75583020e04264bdd14a14e5c"
// synthesis attribute INIT_2A of bigblockD is "256'heb8a9bada32b556a0352bc71f4f635ff1000acb8bb2615026fdee543d4c37db2"
// synthesis attribute INIT_2B of bigblockD is "256'h72d547e9cddb10f3bc2ab1712c32ad51c23a0022dd381fa9d0a8105443eea292"
// synthesis attribute INIT_2C of bigblockD is "256'h3048e1c039d7d21cefc57f8511070a0bc88503ac81bbae7b99b34db6c77c52de"
// synthesis attribute INIT_2D of bigblockD is "256'h2623f94335637969f94ae53849b9d8b4b882f9f35c77c68e664b00c46a84534c"
// synthesis attribute INIT_2E of bigblockD is "256'h99dc8db602a4af8819327d88d72db9fc5f33b65fb6490ee6e26cf31511b9ce11"
// synthesis attribute INIT_2F of bigblockD is "256'h000010027002f574ac1b69daf2187823189959c82fee747aca04587940baf4e6"
// synthesis attribute INIT_30 of bigblockD is "256'h7ceb6cedd91213022a83d46585b642ea845508267c870616640fc81a30f30311"
// synthesis attribute INIT_31 of bigblockD is "256'h1a9aeec3ebec04ba1fd71ff78113eb8d367111b995ebf18f8f5512a1377b8d18"
// synthesis attribute INIT_32 of bigblockD is "256'h5b9d22e31dc2d1854cdc0330f9007274fffbd8c5c4377b5b1d2ddecee56ee9d5"
// synthesis attribute INIT_33 of bigblockD is "256'h58562358074ba7fdf17f870137a1141964038c6e6875207573261939160d0582"
// synthesis attribute INIT_34 of bigblockD is "256'h93bcdb578383edbd8eaa91b438dc3800321cb3dfc999cc672ea6cfbd6b3caf33"
// synthesis attribute INIT_35 of bigblockD is "256'hb8a403ad120c3d5a5741485012263408226822136e01009d04000300cdc61fe3"
// synthesis attribute INIT_36 of bigblockD is "256'h9bdb5cbb14d3f989709bd9b17aa26465998259414b296d56b62d67be757bb5b9"
// synthesis attribute INIT_37 of bigblockD is "256'h860edc95541299b9dca94e878d45b530d35f8bdc93a300332db0dbbe46b40056"
// synthesis attribute INIT_38 of bigblockD is "256'hec2e73b11a4d72496000d8b08cc5412fc6579b6afb3e7a35c913854a919cde5a"
// synthesis attribute INIT_39 of bigblockD is "256'ha887224641e19585001414093090d41c445540ac19f29e85f47f965dd33d0d39"
// synthesis attribute INIT_3A of bigblockD is "256'hfcc13bb45b318bfe95a365876425ad7d48dd96496da1d480dd219223c2d22181"
// synthesis attribute INIT_3B of bigblockD is "256'h9174f371d194dd1027c8bab822dbd58e5fbca82884377751b382405d5b34587e"
// synthesis attribute INIT_3C of bigblockD is "256'h29835c0e18665b7721631e4a91885edb0371fc807274fffb52927cc3be96a501"
// synthesis attribute INIT_3D of bigblockD is "256'ha8522491000716e52d902ee2bb9e7dfcea5be58f8830e814066d2051ac796f84"
// synthesis attribute INIT_3E of bigblockD is "256'h366406ac00023000c34791606cda4a36f127f68e724932b30f53c889e607674c"
// synthesis attribute INIT_3F of bigblockD is "256'ha1e133f85b0b52071d47ce3d525c845c3951b421d608314982a138491440f473"
// synthesis attribute INIT_00 of bigblockE is "256'ha841e5057a735f62596db0a4e4d4887a30cf6a0cf9c100c96e71d8c2c0c94f3c"
// synthesis attribute INIT_01 of bigblockE is "256'hffe2ffffffffffffffffffff9fff4136f6d1b7a8eb675beff6e87f576c67b6bc"
// synthesis attribute INIT_02 of bigblockE is "256'h840006d1547f064f995504e7965f8c43562df2cb0484c542531daa4d24711007"
// synthesis attribute INIT_03 of bigblockE is "256'h0b4384a9988ab1a460c1a20fa43014d429a413a1ba331a95101f9a4ea1380921"
// synthesis attribute INIT_04 of bigblockE is "256'hb6137f8f0e92df3e655a71217b86076f5f8d90359314430125f42a268f544aa0"
// synthesis attribute INIT_05 of bigblockE is "256'h1399bdbc46c439248a5dcbf9fcb8571d09487fa4c1fa1219ef97ed440b511d31"
// synthesis attribute INIT_06 of bigblockE is "256'h807a1c586b465d0f0e4c05229b571ca22f8ac9875a5a038ffd007074fffb30de"
// synthesis attribute INIT_07 of bigblockE is "256'h4dadc5aae41d57704d4739241004bda8dbe777ad5c08a4f62a208a485c908aed"
// synthesis attribute INIT_08 of bigblockE is "256'h56c90fe1104ef61002e2100000645c62f0a1e544ee1c3144bb411a4bd8d34c93"
// synthesis attribute INIT_09 of bigblockE is "256'h837e5a99df6e1393ff40ac2c55aec86776146874c9864e6fb0c71de2761ae263"
// synthesis attribute INIT_0A of bigblockE is "256'h89f7fa2aa61bbb3616206fe851bbf6a1e654e07e596190bfaf15b22efdbeccbf"
// synthesis attribute INIT_0B of bigblockE is "256'ha3349548c281e0ea6e1e931b02090d78ab7b6dc29226f674fd8fa805e15e67a4"
// synthesis attribute INIT_0C of bigblockE is "256'h240045282a7c91e382f2b09a83047c234163b2c49e2a2b8e5f316c661a971ad0"
// synthesis attribute INIT_0D of bigblockE is "256'h7feb8f1dff997c6f345fa7b255b9477b3d4807de990688acb86000b004b04000"
// synthesis attribute INIT_0E of bigblockE is "256'h30d65f1ac235287ae621866e3628fad91707dfdae6492fb80ba30cfd86a7f68d"
// synthesis attribute INIT_0F of bigblockE is "256'h74fffb72d2ff0c817af837746f793a5fb4e80a1ee6ab51d3764a81c91df9a2fe"
// synthesis attribute INIT_10 of bigblockE is "256'he0e2960c2d1c800b71a0462521684df9230e4705e29b201e883dda393b438003"
// synthesis attribute INIT_11 of bigblockE is "256'hc374190f4b7f08d6f36b567870cc34f96b2b094c21c5ba0a1b7f0cc9ef41b4b1"
// synthesis attribute INIT_12 of bigblockE is "256'h55bf705ae4afedf1613a322d802340302100de59981d75614d6d9fb9f7389687"
// synthesis attribute INIT_13 of bigblockE is "256'h6d16e50ce0a467308b487b8c369b685e931ff2f2655c7de23c1444172acb414b"
// synthesis attribute INIT_14 of bigblockE is "256'hf804eff6fe33c82a8bb2affd0b7f7ff3441c5946116bad0e59b5a1a06933734a"
// synthesis attribute INIT_15 of bigblockE is "256'hf19adad652ee8edbd219ee5d2eba79e5402cec99fb408db8a6637ffc9a72e1b6"
// synthesis attribute INIT_16 of bigblockE is "256'h1281292294460925bb746ae1158ecb580d11d8cd090da016b1306abca156cdf8"
// synthesis attribute INIT_17 of bigblockE is "256'h81827d00c4d093cf847837e321055cf38f4806321a1f2ae6f971b068b0c852e2"
// synthesis attribute INIT_18 of bigblockE is "256'ha8dc3b1b884d73ac12939420fb4761faab054b8a37cff5eed8c148bfe1d3b1bc"
// synthesis attribute INIT_19 of bigblockE is "256'h5b39fd43800274fffb723dff90276862f992ef6fdf49a29466f7fb95e55bb2b7"
// synthesis attribute INIT_1A of bigblockE is "256'he8d1db4c0028215061aa6d8cad92f720462c236d0c19024e6725449ba82d863d"
// synthesis attribute INIT_1B of bigblockE is "256'h0e5b7baeb2f9d83e40ca741f52c76db94e3e4e956b0f930c17f38f6af074a83c"
// synthesis attribute INIT_1C of bigblockE is "256'h2767a053ea2c10e008b31166a29584c817911a820acd144001843e42aa7ce0c8"
// synthesis attribute INIT_1D of bigblockE is "256'ha79b197dda70475bea0f4bde4551c744854f176c2795cd3e369245ae71cf9aa1"
// synthesis attribute INIT_1E of bigblockE is "256'h294f3461e5bb2c9e6a5251c7edd3fe8c1f2ddfd7bf518d164ae653cd45f16177"
// synthesis attribute INIT_1F of bigblockE is "256'h9a6fa4a09188fa56991ce475117d39de3f0b0b1c8e8537ff9c8e0810fffcffff"
// synthesis attribute INIT_20 of bigblockE is "256'h15eab492c1b84906b925030a4000791247fb00b12f4fb28bf281e695aa03a546"
// synthesis attribute INIT_21 of bigblockE is "256'ha834f6dfd907d76b16f4b54622c5ff029343929571d62bf896326d0d7a643268"
// synthesis attribute INIT_22 of bigblockE is "256'hc630717c88adf421c3c495642c71cd348c7180926f635935330b91919263ee6b"
// synthesis attribute INIT_23 of bigblockE is "256'h851b9032e93c5a39b63e000274fefb72daffb7efafdace20b1e972cc5b4f6b3d"
// synthesis attribute INIT_24 of bigblockE is "256'h2ef32c6435bc92278e6d4577995ab12a6d0cb192f6c066200f680bad4bc24324"
// synthesis attribute INIT_25 of bigblockE is "256'h1080f03fd1361247aba5ae2fbba8ef89838ce62459943fd81b8d69c9827281c2"
// synthesis attribute INIT_26 of bigblockE is "256'h1ac118a5519a27a955c65db64b29c789d27258f48e8b10cdf42e9c1f0005b100"
// synthesis attribute INIT_27 of bigblockE is "256'h8cfcc3657e31d974c351bde0fea20f0d52fde177ec33b2a3ffbacf555d09ca72"
// synthesis attribute INIT_28 of bigblockE is "256'h8ede0422459136a55ef206b58c45b6ee5a8a7f76460a25a8112ae59e4c6eeb0f"
// synthesis attribute INIT_29 of bigblockE is "256'h0c56a5e19f4ca2a16185eb6a37311b6b2a490801f5c0d63bd632d0bc49b6f8ed"
// synthesis attribute INIT_2A of bigblockE is "256'hd5bbdcfced5db552ed08bcfaa1ec000096c900046610a4d3bf807e8631f7c9f8"
// synthesis attribute INIT_2B of bigblockE is "256'h9375a357a1b1086056cfe2152bda5042881b254dd172bde1e5cfe1dd935531d2"
// synthesis attribute INIT_2C of bigblockE is "256'hebe8098cd37b70ba3b50169b3af11f55032f0f5051ad1a4cb140f1fa8bf13308"
// synthesis attribute INIT_2D of bigblockE is "256'h4ddda8a66718c4bbf82d2639db39ee4d800274fffb7000ff509332fa0d1a31fd"
// synthesis attribute INIT_2E of bigblockE is "256'h908a50e586c552c988987fdb6627722ff6c0d0556119ed8c6a8a0fe064ad376c"
// synthesis attribute INIT_2F of bigblockE is "256'h0e27000080c0c80cadb0d21e13692aadfcb5a618daf42052a4cc2490e3457638"
// synthesis attribute INIT_30 of bigblockE is "256'hbb91026fde2140e298f9b022966a0c907e436508a3fceae3e181b231ea46ad82"
// synthesis attribute INIT_31 of bigblockE is "256'hab41938fe1b3760965ddac9338533653961430ff979093ed4c3f213819c20ef2"
// synthesis attribute INIT_32 of bigblockE is "256'h8fbbe8a59bbcbd092bea5edf162bd749a37eafbec54b742c87dba6c82e6c2241"
// synthesis attribute INIT_33 of bigblockE is "256'h8c21a385863dad9589b98d2327ec1e456891416324ab36af249280109a9f1473"
// synthesis attribute INIT_34 of bigblockE is "256'h933011bc8e12eb78790da960e6834fc93d1a8e96043d000000014412d1c72327"
// synthesis attribute INIT_35 of bigblockE is "256'hffaa53a512bdd8566a325fa133223484f8e708e5ddbdc0eb86b295f5f94c611e"
// synthesis attribute INIT_36 of bigblockE is "256'h3aaebfe63689274dabf9d0663e9bc287fedf64aacc1b9cb680df34b743e6048b"
// synthesis attribute INIT_37 of bigblockE is "256'ha871a4f46da7f121764d2466bb6a1f822e3a398b4cdb0362ff807274fffbbd5b"
// synthesis attribute INIT_38 of bigblockE is "256'h98c00985b0f68ac86cea3923022e000003b527795914bd53ffff0c699c138aad"
// synthesis attribute INIT_39 of bigblockE is "256'h2c36a29c510a0f10000200001f8089a3147fe89c7722df76823f25bbc3b06bb5"
// synthesis attribute INIT_3A of bigblockE is "256'h77463e70def7b5a2ff9a7ea44c2eb3531d7256d3940d70a2424952a7a7233122"
// synthesis attribute INIT_3B of bigblockE is "256'h2856cd4af5b384b007594772cc03355a4c4f702be29e1352cab35e389b1f66a4"
// synthesis attribute INIT_3C of bigblockE is "256'hfe0cffffffff67ff66729e17bfc76a5b7227e6fad9471ceff5648927ad104d8d"
// synthesis attribute INIT_3D of bigblockE is "256'h60127d88946d674fa52cca7899b934901018fdae1b5a668741d40acada439248"
// synthesis attribute INIT_3E of bigblockE is "256'hfe7056ed161d016962aac462a7e355c58901512c158235c7a979003b0000d003"
// synthesis attribute INIT_3F of bigblockE is "256'hb16275f5dd1ced757d0878c3a65773f8f4ba6c29bfd45669fd8fb68152d2a86c"
// synthesis attribute INIT_00 of bigblockF is "256'h7274fffb77d241324cb931a61c3f5ccb977e8584ab2859c8801ca7c474cd739b"
// synthesis attribute INIT_01 of bigblockF is "256'ha54028908aede88c2cf86946ed73a00c2422cb4720626c5831884cda0349fe80"
// synthesis attribute INIT_02 of bigblockF is "256'h92c28c87f51491c38e990f90132cdd259248d64ceb197f2990f14bee7a8f3adb"
// synthesis attribute INIT_03 of bigblockF is "256'h0582d38485e9d6e227e91fae1f331da9083611040f1ccff8568234c5a6a8b5e4"
// synthesis attribute INIT_04 of bigblockF is "256'h9a23525a770d6dc67262abd2331fa7ed3795f5e46a4151d6958e87f68f18bcd8"
// synthesis attribute INIT_05 of bigblockF is "256'hffe9df675f4e7fea7a4766a3ef42e72da844ecfc994c1b3d8395fcfdd421e88b"
// synthesis attribute INIT_06 of bigblockF is "256'hc558444e0f0b86130bcfa80b014434340e99752836dc010afffeffffffffffff"
// synthesis attribute INIT_07 of bigblockF is "256'hc000a82043d071f7e0e473ad4e12c9bd09e7825d6c7ad0f10f4031226ac3f4ef"
// synthesis attribute INIT_08 of bigblockF is "256'h3c4f1b4b92086bb509c9183f61748e1790ccd1820148e27f52f017478bd7871b"
// synthesis attribute INIT_09 of bigblockF is "256'h37bb688315714567784f448053a9bbad88c7bbfb9dc967414e9e375d0a05fe98"
// synthesis attribute INIT_0A of bigblockF is "256'h47d9035fff807274fffb0a36d001c7a35b3cce35437fdfd1daec15bfb2c9147f"
// synthesis attribute INIT_0B of bigblockF is "256'h10ca2286dc29a030cc148aece0803d4f6726150d1c0d0d28cb3321625628b98d"
// synthesis attribute INIT_0C of bigblockF is "256'h0cd5d46088a6945a18197ba31fa01a7bab02949b88312c664a1a0fda49088076"
// synthesis attribute INIT_0D of bigblockF is "256'h06a153776d7a8141728a625a472309672c3d8446005118084068f6933239b738"
// synthesis attribute INIT_0E of bigblockF is "256'h308477620b567348aad9b6317a54804fa0cc10af7f674030aaacb1d6e72d82c3"
// synthesis attribute INIT_0F of bigblockF is "256'hfcbfef6f3b6ee6eae92a95db3ce0cef4c443ac044b9a413757ce79afe540cd26"
// synthesis attribute INIT_10 of bigblockF is "256'hcdb818a6ed8828d252652648fa4fdd4740bb0cc141e4dfb44e3600010000a5a8"
// synthesis attribute INIT_11 of bigblockF is "256'hb2ff6bcb80560925820065a70947407e5ecb6224a838657871caab813eac9890"
// synthesis attribute INIT_12 of bigblockF is "256'ha1f085d2ea9a36d4414d91688b4cc9f515ad35375bace1e73ccd1cf2d0c90211"
// synthesis attribute INIT_13 of bigblockF is "256'h9ff9ffa83d871325a670677b3d7980f1e134ff99da7dffcb27e33217f4bc14b6"
// synthesis attribute INIT_14 of bigblockF is "256'h34c53c4011eb43d902d7ff807274fffb00044c00007af4e8dfed8b3f2b99bfd0"
// synthesis attribute INIT_15 of bigblockF is "256'hd05fd7cc975d3c0a6eb2071baa298c9293ec40c025b16466c90fa00a24271b23"
// synthesis attribute INIT_16 of bigblockF is "256'h009950e08f0a34de3dff0987d769c290f7624da9a8a7a66ee10e81c3c8eb42fd"
// synthesis attribute INIT_17 of bigblockF is "256'ha1880cd538cbdba0d42d8f0356254647e08a020eb18d01e8804010009130eb45"
// synthesis attribute INIT_18 of bigblockF is "256'h6a57989634c94fa536b59a93e271be8ac6c5659526094c2b01343e7b168ce7ac"
// synthesis attribute INIT_19 of bigblockF is "256'hf7f897f4e9479b3aa9ababd800447729645f40a6b3b08524796d1ef5a04a1dfc"
// synthesis attribute INIT_1A of bigblockF is "256'h36a8a8c35294aca99890934a2a46fa08ffff51ff06cf656ac2ae1f7eae71edec"
// synthesis attribute INIT_1B of bigblockF is "256'h1894d9dc0310203d00002004846be8884097b5b6a626622c0e4836668eb6af76"
// synthesis attribute INIT_1C of bigblockF is "256'he9890f3dcc5426774efa06e0ed5a4b9f4dbbad48074cc08f0e57a6796407a76b"
// synthesis attribute INIT_1D of bigblockF is "256'h5ce66fa987e690d1bcadaab233e0eec584f89b95ffa9ac5aa558ace8b2969cb7"
// synthesis attribute INIT_1E of bigblockF is "256'h7c4a24ad9b3d34c43db0d18a3e5902ceff807074fffb3f82ed7982b7a6b706cc"
// synthesis attribute INIT_1F of bigblockF is "256'h35d69fdf01201722caa59ef70e0f5e55ab85a1f1e8c313ec80cba4516747d8f9"
// synthesis attribute INIT_20 of bigblockF is "256'hbbfc0054000087aa07fa22430a2b8e3f755a4a508b2a7615189024095d8e447c"
// synthesis attribute INIT_21 of bigblockF is "256'ha285b30355ab36341a7055eeb26865a5c374368974ea14ae131df408f9785184"
// synthesis attribute INIT_22 of bigblockF is "256'h35f6281ab1181442a410ed55a3639607c4d9088269b7515a197893d8ea5e526c"
// synthesis attribute INIT_23 of bigblockF is "256'h29ff09c23e860a969166b21e7dc790ee0afe7fc8ebabe4650ed4c5628e2cc590"
// synthesis attribute INIT_24 of bigblockF is "256'h180e502cf48203dc322a18ae5d166a7cd066d43038c11f85e6aa0002f800ffff"
// synthesis attribute INIT_25 of bigblockF is "256'h49185c4501042789a446476cdab60a95000000007283c999d3fd88750cb1912e"
// synthesis attribute INIT_26 of bigblockF is "256'hd3bbc3c548601fb52f981f36075220b27ea1c3cf01f841ef1b0691780129fcbb"
// synthesis attribute INIT_27 of bigblockF is "256'h1517cb7bfc66fffffff8ae1b858b6f8a6fadcebd7ea68effefb421b8ae2aa4cc"
// synthesis attribute INIT_28 of bigblockF is "256'h51e0e7a40d640c65a982273022bbd824e914d9516d4d000374fefb72aeff1e6f"
// synthesis attribute INIT_29 of bigblockF is "256'h1d4bc40c6efaaaa063a1893bae9b003fc2b0e585c1c320390896928eec88788a"
// synthesis attribute INIT_2A of bigblockF is "256'h26e1ae5d809c000000000100499aaa00c277b352aa9365842616c40412048bde"
// synthesis attribute INIT_2B of bigblockF is "256'h2b0be0b650c3b92242c83e0a91312dc6c294c12f4637d063a2b85f098e40bf55"
// synthesis attribute INIT_2C of bigblockF is "256'hbfdbef1f8f129ad25f2f5db9fada9d5c053a6b1d41784fb299087172466442e8"
// synthesis attribute INIT_2D of bigblockF is "256'h3ae5d38bce75a6d8b93e66637175588ff98d3ad2ceb245619aa9323ce44e1e5a"
// synthesis attribute INIT_2E of bigblockF is "256'hfffd1fe37cef1ffcf5ff0c988d8c336c55c5a45ffbb19e9e5abbff9c62f3718d"
// synthesis attribute INIT_2F of bigblockF is "256'hffff81ff70cf3e26f713f4bdffffff5ff3ffebffadef358fa7c6677af37aa969"
// synthesis attribute INIT_30 of bigblockF is "256'h1231c2330f2385a97a8c5da11540561268627f3cc98a2187ecbda285dd22fbf2"
// synthesis attribute INIT_31 of bigblockF is "256'hfb7278ffdb343b528af23f674d9ab138903015ccc6d131b492ab246962f37595"
// synthesis attribute INIT_32 of bigblockF is "256'h98606c1a9288000054c40d610c05c9740930c2bb6828862c58194443800354ff"
// synthesis attribute INIT_33 of bigblockF is "256'hbc1ae63c005ff52c6bad148f6687976dd6ed39e5e090213445500ab3000c01c0"
// synthesis attribute INIT_34 of bigblockF is "256'h3295fb5a14cd7769381ddfccf3ba37cf48e0de362e4998a2707539a8a2806ac3"
// synthesis attribute INIT_35 of bigblockF is "256'hc0575295a14c82c2695342202f90f401da6cff730ecaa1bd926557d2c5208cfe"
// synthesis attribute INIT_36 of bigblockF is "256'h4a3cfbbc9656b706154a8ac50820bf90cd05390b1bb11c0a94457333e3a4e96a"
// synthesis attribute INIT_37 of bigblockF is "256'h1572d07ce636fbb2f88e14551de5e3f98f6f6ca6d2b923145248f18c471ded31"
// synthesis attribute INIT_38 of bigblockF is "256'he11d8caadd1593ddb12dbbbb05bff4aa6a86fa7886dd5a5bbb3bd35d1591dc0b"
// synthesis attribute INIT_39 of bigblockF is "256'hc7682fd2ffc28d7fa7a12927afc2eee5ffce977fa1a46e0331974b25578d97cf"
// synthesis attribute INIT_3A of bigblockF is "256'h402a1442280fc24c3f8abb525538ccaae500d32afff9ffff90014de90cfce54e"
// synthesis attribute INIT_3B of bigblockF is "256'h4164800574fffb72afff8386258852604a5c413c08bc2e3a8a9ae0ef98023f2d"
// synthesis attribute INIT_3C of bigblockF is "256'he22d019900121ec02b8b078f0001399c915c1cb9bc00e2c743ca00413de05736"
// synthesis attribute INIT_3D of bigblockF is "256'h0919f7ac19660634d2852720015c925212224204e13a194b62b250cd0a042c8d"
// synthesis attribute INIT_3E of bigblockF is "256'he1e62eb841e3977b4270ec725235411d8ed4810b5b9a87c8300750ea108aa056"
// synthesis attribute INIT_3F of bigblockF is "256'h79976dc863d6e356fddf7d75553277cd577c476f70dc7dd7495518646bfb20f4"
// synthesis attribute INIT_00 of bigblock10 is "256'h46f92492a6b7bc0070c5e9adc045fe13e63d2e78dc9fab32cc4c0f1775c78ebc"
// synthesis attribute INIT_01 of bigblock10 is "256'hb05ba6d0bbd8c51db7aee84200c2748005fd6846520aa910a25893525b68f252"
// synthesis attribute INIT_02 of bigblock10 is "256'h4d315253ecee1ce29462978f25f0571269b4f2dd9cb7e044d5635a7dfbd9ca15"
// synthesis attribute INIT_03 of bigblock10 is "256'h0f5a19f5ab33e6eb7ed7367e00f731ef5db32291bcd330cde2c16e2d8ab34001"
// synthesis attribute INIT_04 of bigblock10 is "256'h4f3efc12a4a61b6d85134c02f59e7e57f31d5d178b1a1b2d4d5550bb2e2ef7ff"
// synthesis attribute INIT_05 of bigblock10 is "256'h0a153d00dde75e5000037482fb7052ff171b00154ac027236800b0930ce9abe4"
// synthesis attribute INIT_06 of bigblock10 is "256'h3bbae443ca5b6aa5ad5908bf008c6ee84905d8e8260c25770cdd8c00bae0221b"
// synthesis attribute INIT_07 of bigblock10 is "256'h878786853239e466da0cdcb1420c645dae826ed14e3e54ac5084f2bb2cb596b3"
// synthesis attribute INIT_08 of bigblock10 is "256'hb420223c98f5eb1f34c33b79e7b697b48569b3b9d50c85fdca88b9be46b028ad"
// synthesis attribute INIT_09 of bigblock10 is "256'ha32f5088d9ed7d00db4a51b6a491003047489dfe9aaa9953ee7b25a339b41801"
// synthesis attribute INIT_0A of bigblock10 is "256'h686a8edb1124f52a7980e236a3a9b5679c0e0a92711006860e479e80b4784337"
// synthesis attribute INIT_0B of bigblock10 is "256'h5d5adc6a311669bef3b663320597bbd04a6c3528f645e392106e588ba87e1db4"
// synthesis attribute INIT_0C of bigblock10 is "256'h4b1db3a1851730d4ab14fcdcec3c1f5ef3769e1cfa7522f3e71796756f24a564"
// synthesis attribute INIT_0D of bigblock10 is "256'h1e263a304f3ed43b1132c9ac7f26d2417236486302559ab6826cdf336ac3fb19"
// synthesis attribute INIT_0E of bigblock10 is "256'h9da1575f9ec6e85da9b926090ae83b14ccd5c376d09439e8000949a0326a1640"
// synthesis attribute INIT_0F of bigblock10 is "256'h000c00221bbd15021dbae185455d03278f807274fffb9bb33ec219e8efd18494"
// synthesis attribute INIT_10 of bigblock10 is "256'h526a6630974a4a3678ad5a8a4a11364138590d80f413086ec85e147877e69535"
// synthesis attribute INIT_11 of bigblock10 is "256'he5fcbdbec77763280d74ad9d6e0e84b674a16a93332e2b65ae74a7e1936a32d5"
// synthesis attribute INIT_12 of bigblock10 is "256'h5880a800c006852b1f42944a2c0e6e0523941b6d1049011c5997b2facc611ecf"
// synthesis attribute INIT_13 of bigblock10 is "256'hd4419fc9ff88c0f7b89e52bace7c90ffa073901fd0be3d50865c8ab8a89c070b"
// synthesis attribute INIT_14 of bigblock10 is "256'h94d67d4555c30cd4d44f1fcac3b6e07c3b3d534b3bf94afe22d9676f82bce9bf"
// synthesis attribute INIT_15 of bigblock10 is "256'h0c28e82a5bfb4d9b85c0ed7917512db60c47baa307d8f72a55189a470447294a"
// synthesis attribute INIT_16 of bigblock10 is "256'h9c6d20226d860541293a49e60611e78450b6a463236d2949010950094e1b7040"
// synthesis attribute INIT_17 of bigblock10 is "256'hb728798223b15f919d3a2ac9c2b57c14f5384e0c4d31ac09cb5d116a0019a000"
// synthesis attribute INIT_18 of bigblock10 is "256'h51e3a29d63149c81acda9a078cab50c109ea53d1c5119e3d8e06bd984c6017d0"
// synthesis attribute INIT_19 of bigblock10 is "256'h24b671864d19180d00261b8a124115a269874cdc03189f807274fffb13b4cef9"
// synthesis attribute INIT_1A of bigblock10 is "256'hf6d733bb0f95a2e9f341d16cdcdfb5225b617a2a99d5f35d88203400896ee05d"
// synthesis attribute INIT_1B of bigblock10 is "256'h9cc18bf777f000bddc3f0e114e189fa48e3619241b61e00366644ae7da1480fc"
// synthesis attribute INIT_1C of bigblock10 is "256'h2b356cf69fa1044a8a81547ab51960f09eb05a14b92680125380c1b84e00cdec"
// synthesis attribute INIT_1D of bigblock10 is "256'h1d2bb4970c6e6d67a056f04f4514ed0c6aa16e198b0d0f859d0375682148dbaa"
// synthesis attribute INIT_1E of bigblock10 is "256'h19813c792cf86b59dc1050e3c3406ca96df02a3f04ab2b693ab16a8bb34d76fb"
// synthesis attribute INIT_1F of bigblock10 is "256'h014b94005c540a01195fbc6b3df787fd6f6e71f5295f20c26da94924c859a801"
// synthesis attribute INIT_20 of bigblock10 is "256'hca98de93e384f7d2dd09a88bc87680c73fc4d1c4816e86c12176440d32a45981"
// synthesis attribute INIT_21 of bigblock10 is "256'hc6759b3b3da97fec83a63d386516c83a5e5d9c295c282adefe06f4f6be1fe21d"
// synthesis attribute INIT_22 of bigblock10 is "256'hfffb0104f81844a9b241d43b67088e160739f4b36da876a64f31d2d5517f35f9"
// synthesis attribute INIT_23 of bigblock10 is "256'h2801096e00609c5671a4c4d90a0b00685b8d1a82155a69874a5c0343af007274"
// synthesis attribute INIT_24 of bigblock10 is "256'hca1456e22ad37327eeb8e0d911b56d1df4223c13324a836745066d6ba31b1848"
// synthesis attribute INIT_25 of bigblock10 is "256'he7dcd4e01e55ef50068b0fefbac99281feeecdb0f192c0905c60028500000220"
// synthesis attribute INIT_26 of bigblock10 is "256'h3ff9658f6e3c3ec3b761e271407ef8d61cad6ff02c59e29ac51fe384bad50202"
// synthesis attribute INIT_27 of bigblock10 is "256'ha2e0bb415d62604d614e78ee9672ace94dac57e38ed4eeb93cece7df088e8569"
// synthesis attribute INIT_28 of bigblock10 is "256'h9d3b1deecc632669054c020014b08d55c78f1fc541298471b45ddc8d00482040"
// synthesis attribute INIT_29 of bigblock10 is "256'h57abfdb8bb918339519e97b10d7dea87897f95fed08e6bd61c5c506d37c5a4d9"
// synthesis attribute INIT_2A of bigblock10 is "256'h8ab90ee465904815f6f9efd02b21019c5851405df50528adf63c001ac6cc6926"
// synthesis attribute INIT_2B of bigblock10 is "256'h105dbe03b6262ee978f746842465e48d08b81404d4605da5cacc2357e24f2a2a"
// synthesis attribute INIT_2C of bigblock10 is "256'h030dbd807074fffb78581dea8a66af3128368c4518a3f2d5c2f9005609402ca2"
// synthesis attribute INIT_2D of bigblock10 is "256'h29ee9ea38c003400852ee046a051714411352c0c04623b8a2044436850c942dc"
// synthesis attribute INIT_2E of bigblock10 is "256'h8f258850c3a163175491fe20f1525233d1950d2ca26990f226abcd118f09fc3e"
// synthesis attribute INIT_2F of bigblock10 is "256'h91d544b399c855f5b436a0d972ada54166ec7a96bd6f0872704cdbe6c32c5cc6"
// synthesis attribute INIT_30 of bigblock10 is "256'hcddd00271432112bd005a1316915b8db806961421e014f17a8c2dde872e53edf"
// synthesis attribute INIT_31 of bigblock10 is "256'hc9330452cb2a94d308904a2b002548025400c2000a44e452b1743f5041ee0590"
// synthesis attribute INIT_32 of bigblock10 is "256'h471530b5a77f8d8f2e3e1fe6c033e16c8c23ad4e87b96ea59b1536684a6fad36"
// synthesis attribute INIT_33 of bigblock10 is "256'h0b78c895810ce500a4cfa247bd060a11561f2a4219bfaa8047fc2e37ea1f1a4e"
// synthesis attribute INIT_34 of bigblock10 is "256'h161f815d5fb11a6992370002c03c0519a32a8a1fba0764474cc40605d9461a90"
// synthesis attribute INIT_35 of bigblock10 is "256'h30a78bab32ad8fc6211c4e3db05838b02990400101a448452c80ab18e940b6c2"
// synthesis attribute INIT_36 of bigblock10 is "256'h081225175cd1d33e000274cefb722aff80b96d5aa8bb077dd2ebe39ee6222c6b"
// synthesis attribute INIT_37 of bigblock10 is "256'hf1d83cd194cc8b80f30631f60194ee74888c51e0a62075734d19490c9d00c16b"
// synthesis attribute INIT_38 of bigblock10 is "256'h32b3846f31ce1cd4e933455aa2189c63fd67b320733fc1246182883f453045d3"
// synthesis attribute INIT_39 of bigblock10 is "256'h9d0ce77a692426db112ea70322a819c607e5322953fb6391d9aa636d7b4c57b2"
// synthesis attribute INIT_3A of bigblock10 is "256'h5a98fbdb4c8f95637137e08a9dd1496901431200000a240f9e612b24e935a0f9"
// synthesis attribute INIT_3B of bigblock10 is "256'h1725cf5f48440ba6ffec2b6684a7d7af14b6db1e5c48bc7d19665ef058cbfdd4"
// synthesis attribute INIT_3C of bigblock10 is "256'hfe15c49f4eea67b79482bb8991c1f7a99802ef504d77edb83065e35e98c9aee8"
// synthesis attribute INIT_3D of bigblock10 is "256'hb68b148d0040bc38e982b243ca84af047ff8d78cf05d865a8a49f8bf8dff6ffe"
// synthesis attribute INIT_3E of bigblock10 is "256'h97104020c0483c1e0f036b8c844750f3d62b3de98f43d0a6adfad62549330b2d"
// synthesis attribute INIT_3F of bigblock10 is "256'h32b7f0ab6ac7b4287a5d26e2ee333d51433476b5a5fd69931ee82e1bd3388648"
// synthesis attribute INIT_00 of bigblock11 is "256'hc5307d0c21abd0158b1cdbe92a33000374ddfb72adff600dc774d9d4b246e367"
// synthesis attribute INIT_01 of bigblock11 is "256'h6fad37f462865ffb4234ae9a6727bf5da8271494ade85006b608a62c6d6f0d35"
// synthesis attribute INIT_02 of bigblock11 is "256'h4200558975bddd5dbff5295ab3fe5b41aad2f7fe5319fd6ff8d7dd8fa2f91d0b"
// synthesis attribute INIT_03 of bigblock11 is "256'hac3448b9d17b00200020004092896c213154fe7d02f5bb0a9843ffd202773200"
// synthesis attribute INIT_04 of bigblock11 is "256'h53e7cea652b3d971d4e0be1d61dca235d2a8449ca95666b49cf10891cc242e96"
// synthesis attribute INIT_05 of bigblock11 is "256'he54fc107ee5ac95f2049c8ef1d45fa72301fe9d7aba9cf013745efdc0489b69f"
// synthesis attribute INIT_06 of bigblock11 is "256'ha7b199d35ad472a385852d5ce9a3b6aaac8e335ddfd43a908f59b6ea17fad8d4"
// synthesis attribute INIT_07 of bigblock11 is "256'h7e14a21383379ae459be425384a99a89ba05927449260b1340007c04aea2746e"
// synthesis attribute INIT_08 of bigblock11 is "256'hfb33b6a2e9154a9cfbaa959ecaa9aa10c61e4520fe4cb3dc4bda00040000d802"
// synthesis attribute INIT_09 of bigblock11 is "256'h98d54a48296b4d74b110d950318b877ef397ad71ce3c65c1311769acda92545c"
// synthesis attribute INIT_0A of bigblock11 is "256'h47a0f9670c48251e3a0502bb2220e92ed9d17e33000374ecfb7201ffe425b75f"
// synthesis attribute INIT_0B of bigblock11 is "256'h84f52fff8f9e5afff8e7e36f56ea2cc506e6b88ad6aa9023160c6cf05406b888"
// synthesis attribute INIT_0C of bigblock11 is "256'h846edb608f506ab10a750201c915b7d96a88b4b7170c194e5e6aa88beacefe5e"
// synthesis attribute INIT_0D of bigblock11 is "256'h218f59528d25246bc16588f518b800000000c00002001c07a360c6525eaa0feb"
// synthesis attribute INIT_0E of bigblock11 is "256'ha2c87189d7d6926862d362b944bd57b771b0f1734d9ae1e36da61b6c89445d66"
// synthesis attribute INIT_0F of bigblock11 is "256'hf2fa020e846a5afbb9937e2b61b3c288d4540f3c851a37ba7b6e2facf6324cf5"
// synthesis attribute INIT_10 of bigblock11 is "256'h5557000d0d00a3f015cb6998e080b6f987010b5a61a5659627712b6a5f443a97"
// synthesis attribute INIT_11 of bigblock11 is "256'ha4f116cf32db02ab0000008005088ba8540e0517f3e62f7106936289c3142492"
// synthesis attribute INIT_12 of bigblock11 is "256'h4cf50966aadbaf1e1e3da4884c7ff97f82b61ba1149b8523914b07ea41402e5b"
// synthesis attribute INIT_13 of bigblock11 is "256'h0aff59339f5c723760f5902c462ace3e9c82baa371931a87faa1723acbe03f30"
// synthesis attribute INIT_14 of bigblock11 is "256'h6be45c050b808c3d255f0dede908fd05e1aa301beb1657e1865e800374f3fb70"
// synthesis attribute INIT_15 of bigblock11 is "256'h5efbbc16f8629dfcfbff054fa8b93cb176a13647bf09925ff27f57c399e565b0"
// synthesis attribute INIT_16 of bigblock11 is "256'h068700002000dcbaa42d10de7a4c0685cc9362ee10d5a0ccbaa800aea000e100"
// synthesis attribute INIT_17 of bigblock11 is "256'h89750623bc54fa85e50f3c53d31b7198304755a1595d68fe050dd2e1f1c1ebe3"
// synthesis attribute INIT_18 of bigblock11 is "256'h57344c91f62fa1fc0c7a85473ab243162767ad5db6d25f74e687ac89d11a0283"
// synthesis attribute INIT_19 of bigblock11 is "256'hb2366ea7c2567001e5b12353e21e022a2a5d40b09d978b81b8f956672ee28162"
// synthesis attribute INIT_1A of bigblock11 is "256'h9b68efcd93a23b0233bb0430814ba0a42aae555f0015fe00ffff88ff60f3e38e"
// synthesis attribute INIT_1B of bigblock11 is "256'h97bdd76b17506e92dedac1bcedae4ecc69e2b7ae1a90a32ba7302ab000001c00"
// synthesis attribute INIT_1C of bigblock11 is "256'h032ea69973b75afdbf34ac7352ade2a63372b87df0c10b65305dfa8d888034c0"
// synthesis attribute INIT_1D of bigblock11 is "256'h0374f4807274fffb721b2a370a6baf354f652f9d532ba6153c15cbae9142d3eb"
// synthesis attribute INIT_1E of bigblock11 is "256'h2f88f5729888303786ace863b0ab61a76cc9160d05e67b0c184116a869e843d8"
// synthesis attribute INIT_1F of bigblock11 is "256'h7f18a06ad3001d47c5860e484db5b513000121a024797318481d57fe332f93f1"
// synthesis attribute INIT_20 of bigblock11 is "256'h7b5298ea93c4930342cbdfc6602590993c1550dc0000db00ad77b10f945e586e"
// synthesis attribute INIT_21 of bigblock11 is "256'hbca112328a208bc959a112699128a362f939e9607522d10b779cbbbe4d7c2989"
// synthesis attribute INIT_22 of bigblock11 is "256'h3abc8e6a472c0f7607f62c914c5106b0b431e42d64830e3cb7cfd649ca661417"
// synthesis attribute INIT_23 of bigblock11 is "256'hfeaa000bff01ffffffff3e8f6d4389c0c9b90a2dd097194a7a0e141b56fd16d5"
// synthesis attribute INIT_24 of bigblock11 is "256'h2843984d91b3006000002e344504457b78c0a142c66d60bf164261e98b0f84d0"
// synthesis attribute INIT_25 of bigblock11 is "256'h281d142801f88f027119f28e430366881708c3b0420fe4992cce85a0b98e21c4"
// synthesis attribute INIT_26 of bigblock11 is "256'h5472d69580bce8e2e435ad74db089195c93c90f8a03c3a22e2ac41908c090ba4"
// synthesis attribute INIT_27 of bigblock11 is "256'h42f839ec34d70377fa007274fffb78ff6e3dabee857f29f995fda2cae5260e3c"
// synthesis attribute INIT_28 of bigblock11 is "256'ha451f0356746e5a8bfffb0c8a86786abe06eb0af5c671127320d1969aae91801"
// synthesis attribute INIT_29 of bigblock11 is "256'h8b0d4f4348ef4b628d3f75587484d2dfbecab9a88a49322400009000d2ec5fe3"
// synthesis attribute INIT_2A of bigblock11 is "256'h3f8695567e2b59228fa5d7436758994c6c41615b6247042408000000bc04a71a"
// synthesis attribute INIT_2B of bigblock11 is "256'h0e3efdb7da36ef8d5e90ad7b46dfd5a44df73b790aa8d79bf597a6e6a531bb5d"
// synthesis attribute INIT_2C of bigblock11 is "256'h6ffb8c7b2ff31f1156c9be257a3f1b8bb7ffee14111e6397c9314dc6723427b2"
// synthesis attribute INIT_2D of bigblock11 is "256'h0bbb4fe17aed2e5063deff5de77f6a67fff7d7ffdff79b75d2f6bbfba7d6df54"
// synthesis attribute INIT_2E of bigblock11 is "256'ha042085a4b1d797910b5b09d6cc339d0c272233829575478a555c0aa4abfcdb4"
// synthesis attribute INIT_2F of bigblock11 is "256'h54a378442583a39158e385729944ce0710f34a2c89a00190884750ca08a07331"
// synthesis attribute INIT_30 of bigblock11 is "256'h716d058ea1e3c30453880ca69954c42c1672c6f227d20b48cb83343487214489"
// synthesis attribute INIT_31 of bigblock11 is "256'h0d2caad91ae115b899e945d60390ff807274fffbfce64e54f3499c8b697d0b34"
// synthesis attribute INIT_32 of bigblock11 is "256'hfd693e6495cdd42bcc53b3babe76baab6000769e86ab2079f4005a74590f040d"
// synthesis attribute INIT_33 of bigblock11 is "256'h9e547128d47c4d84a5ab16f22a16b85ac51313d26784970abfa00d21b2c95f57"
// synthesis attribute INIT_34 of bigblock11 is "256'h5c81542f9f30b6345a1394fbedada8a6ce1e0b278eceda77c1f7a8bc4978beae"
// synthesis attribute INIT_35 of bigblock11 is "256'h12712e4216a3427118e69c6e166355552aa919d0439bdffeab71ffb37ef79d3d"
// synthesis attribute INIT_36 of bigblock11 is "256'h17d5e832a88a2c854e9188d963fa200cd07342d146253c0e213e428e5d9d0620"
// synthesis attribute INIT_37 of bigblock11 is "256'h8ea46f86f3610000534c00c038c3b2ac1e5fa4465a8d3c98e7d32ad350854a41"
// synthesis attribute INIT_38 of bigblock11 is "256'hde0a6711c5518f97072258e124311d428f23340837521fdf1e925116c8909d2a"
// synthesis attribute INIT_39 of bigblock11 is "256'hb3fcf1b6eb8fb97b6d7f78e26620e6ee1bb8ef6b1491cd4f3067f86676ef10f9"
// synthesis attribute INIT_3A of bigblock11 is "256'h5354ffaac16baffd971f139ce3c65533936d36d6ff2da3fed2d049d5cc73cdc7"
// synthesis attribute INIT_3B of bigblock11 is "256'h5a18050f0011c7a4cad23d23e0009e3d4dd6040aff807054fffb4f345290ca74"
// synthesis attribute INIT_3C of bigblock11 is "256'h5fd903c4e47a0b3b5e3b4f27000084000b80b8bd7c52f0004b1e0f2b091af600"
// synthesis attribute INIT_3D of bigblock11 is "256'h9852bc9ee5f791df24c0bc84a1ffa786c9943825a7b6f47e07b2b0a9787c0865"
// synthesis attribute INIT_3E of bigblock11 is "256'h21a1a0847830dbbc3347dbc44e2e605708691031569806280d66d042fbec18d0"
// synthesis attribute INIT_3F of bigblock11 is "256'hd755000d36aca7170e3e2848ab98dd6083e1db10d506b024acffeeff3deeaed3"
// synthesis attribute INIT_00 of bigblock12 is "256'hd89799f70aa88e413c0a90257084125b1b9288414299b1cc209a42c952a71f27"
// synthesis attribute INIT_01 of bigblock12 is "256'h81960a399a88a838369d360a931c27c133da4c72d758477b8eab7b2f484d9ff1"
// synthesis attribute INIT_02 of bigblock12 is "256'h7f45ffb9b5975fc2b19e52fe217917ffdb920736867d52557ce3a9335bfaa15e"
// synthesis attribute INIT_03 of bigblock12 is "256'h9a4949c402dbf8311dc76066b28800c08b2009c3b8e92f7c919c6f1a2a5e7553"
// synthesis attribute INIT_04 of bigblock12 is "256'h56ffe2a856e0b50d503e29d30003cb0a13b5ddb0d2899d5c7809dbce39d92099"
// synthesis attribute INIT_05 of bigblock12 is "256'hada45085d060232c236d4d79000066e3812b081119005b672d56800354c3fb72"
// synthesis attribute INIT_06 of bigblock12 is "256'h3098c9b2696ab83b8bdf1e0bde7465e52d8c7bdfde87f1b08548b4ad8151608d"
// synthesis attribute INIT_07 of bigblock12 is "256'hf7776df36c99e9878fd841120fff523d631595e836995149d456a08c123b758a"
// synthesis attribute INIT_08 of bigblock12 is "256'hd9328a12f540862574a87ee774883eb2c9ac2522f62575815cde9d4ff3f35b76"
// synthesis attribute INIT_09 of bigblock12 is "256'hc5db3b09e5ba3cb08a3500397088a79a2901771db667f2c695d6dcd0491f371b"
// synthesis attribute INIT_0A of bigblock12 is "256'hdb706aaaaec521997fd62c18aff6fa924110548e46b89d5b1225ab3f12285006"
// synthesis attribute INIT_0B of bigblock12 is "256'hbab98f4e516e5918d95c9eccfa5275ac76311b7ee6b5626aca2fc42eb1828b6a"
// synthesis attribute INIT_0C of bigblock12 is "256'h1782c079d42a71b6451b5a29fc022fd9870eea358c9d9d5d969acd764a8a9edb"
// synthesis attribute INIT_0D of bigblock12 is "256'h1202b51107b1cadff14985c73937cba4b0fcd1890c2c6000438b8042f46a4109"
// synthesis attribute INIT_0E of bigblock12 is "256'h000374d3fb7257ff21fe88de11c2f894ff26896780df2604e0016bacbc5d2eed"
// synthesis attribute INIT_0F of bigblock12 is "256'ha69e00b31018aeb44f05d568879c05754d392602ad00e16b2214881ddd694d5f"
// synthesis attribute INIT_10 of bigblock12 is "256'h3ca1b58ef1c1fddbe5b1fc488ff71d93a7420d917eac82667624cecb94e9c06a"
// synthesis attribute INIT_11 of bigblock12 is "256'had66ed8444f6004f34b9d8581af772478284700819cdc5dc976373083dab1a57"
// synthesis attribute INIT_12 of bigblock12 is "256'hc9b7b3eb235d62cdb324d0c898b14a61b40095a5400a555e141a0c948a2efc9e"
// synthesis attribute INIT_13 of bigblock12 is "256'h377058450e34e624c71e59ee942868846615a694a9e98963331122563185a7c8"
// synthesis attribute INIT_14 of bigblock12 is "256'hbf25d4d3febb6a8ff08cb66fd884de4fcc44d57fe8a7a54f400c77e7562be1c7"
// synthesis attribute INIT_15 of bigblock12 is "256'h0e20be776c9685e1b50bfb6b2ddad90866b9eec95fff48954422838fd4969dec"
// synthesis attribute INIT_16 of bigblock12 is "256'h600fc32837b4bfea194bd203d95415903227e20351ec001898c073365bab2ace"
// synthesis attribute INIT_17 of bigblock12 is "256'h20fa5b10f0cf93d9cee00491a71fab6db255404cf06c8570acb29c44e3e09ab5"
// synthesis attribute INIT_18 of bigblock12 is "256'h862ddde11e5b000374e0fb7215ff7ec6a9ba02c2edd11a3ee0a1dd1031f91af9"
// synthesis attribute INIT_19 of bigblock12 is "256'h612ee37f1f576fce415f231e2ee87a0c7a60449817774c810300bd00c12b2a11"
// synthesis attribute INIT_1A of bigblock12 is "256'h3070d4ce2dfbc49d56629348b5631c6d2aa70223040363b30c1f6b7522e3c9e8"
// synthesis attribute INIT_1B of bigblock12 is "256'hc7373bc6fb0127b1d82c25d6240000198c52916aede2105df18d1b53d5b78016"
// synthesis attribute INIT_1C of bigblock12 is "256'h10ed89b4d8a41f38a298fb913886bd14647841147909302ddd63ee6f737284e0"
// synthesis attribute INIT_1D of bigblock12 is "256'hbfadd91fdf31a55868e6f9d476b75960f43db491839709c23698396efa2f72ac"
// synthesis attribute INIT_1E of bigblock12 is "256'h218c6ba5f3ce8db5049c4480101a172471e52a379d73010035ea35d57fea87d5"
// synthesis attribute INIT_1F of bigblock12 is "256'hc40e7a70472c048722002848b6683d6bbd15eadd1b48bef980a6b3e2586eddd0"
// synthesis attribute INIT_20 of bigblock12 is "256'h74c67cefe6b1ad0dbebe6d5b2c9afbde154aac6ceddb296b29566155c6072349"
// synthesis attribute INIT_21 of bigblock12 is "256'hf3bbbac656fe6f4063585ab07b5c27d585aeac7253158bd3d30ca96ab61c22c7"
// synthesis attribute INIT_22 of bigblock12 is "256'hb90982cb121c23165dd1df49000274effb7052ff9894a32a4377b554169a55ce"
// synthesis attribute INIT_23 of bigblock12 is "256'h4eb3d487dabf931aa7e24fe766c3100900a0eee88a8dbe20449c25774ca12390"
// synthesis attribute INIT_24 of bigblock12 is "256'h424d9a54c9f2853d1e315ae2a1906ecefb8a19c1372dd3596e83dfff8410bf88"
// synthesis attribute INIT_25 of bigblock12 is "256'h129786a9b039452df9bdc9ea13960698edc291a13af16116770e2859a04e4517"
// synthesis attribute INIT_26 of bigblock12 is "256'ha1bf5c95672218f11b3adffa9b5e20e9753c440a39c1ca49bd124f3dfd5a4b2a"
// synthesis attribute INIT_27 of bigblock12 is "256'hfffffffffffff57ffa9ddf2b4fa14c6eb72ffe56cb7f4115e3fd925e12c79180"
// synthesis attribute INIT_28 of bigblock12 is "256'h4d43a044cf3606133dfed67771b604008000ffffffffffffffffffffffffffff"
// synthesis attribute INIT_29 of bigblock12 is "256'h0ed18a1d7d278caaac35009f790808629eefa8805e1581d2841f6c0f7e69d3e6"
// synthesis attribute INIT_2A of bigblock12 is "256'h637f9b6e721c33bdca2e72eefb1ef55896cc2518d2f8f62ed2239b7c0b953e7c"
// synthesis attribute INIT_2B of bigblock12 is "256'ha9bc0a5ff485dbdfcd5b5c1b32eac4e99db7656d171df5bcac7df02486724252"
// synthesis attribute INIT_2C of bigblock12 is "256'h71265541640d18287b871ee32db0518848dc032ef9807274fffbfd1a2a68ca43"
// synthesis attribute INIT_2D of bigblock12 is "256'h1c1c61b62296bf39e46d4400ead44feb1bbf5bf429bd8cb918240ceea07f3cf3"
// synthesis attribute INIT_2E of bigblock12 is "256'h285a15400000802689005f96451abcab28f33847435ccad9fe0feb108fdfb82c"
// synthesis attribute INIT_2F of bigblock12 is "256'h121938cd6b25908a558a27e1e0153d83028b76496a300e36f34668a90f174814"
// synthesis attribute INIT_30 of bigblock12 is "256'h31186ccd2775a0f4fdc63291b67f812438eaa223bca4f3f7c0b9a6a58d57b150"
// synthesis attribute INIT_31 of bigblock12 is "256'h9fffbfe22d7e522c3d7495fa27db35558e86fab27d91232a634556cdaee5a0eb"
// synthesis attribute INIT_32 of bigblock12 is "256'he41069ed25880c722b149ef7c53513552caee45935a0dbee2e460088fffeffff"
// synthesis attribute INIT_33 of bigblock12 is "256'h1c02bd9aec30e29bda5c1599ba2feefa9588dafb0eba1d6484000505d47067c7"
// synthesis attribute INIT_34 of bigblock12 is "256'h4364ab11ecb1b9ba9bf87553deb19961f6edbd324a31719ddd3dac6c78e967d7"
// synthesis attribute INIT_35 of bigblock12 is "256'h5bf4542fbd59f433c70dcb6e91aaa063c3c03f76a531077676ccb216ba4c6147"
// synthesis attribute INIT_36 of bigblock12 is "256'h0ded00892c5e6a46b523824b19833b5a25031470898941da0361fd007274fffb"
// synthesis attribute INIT_37 of bigblock12 is "256'h3bd6b00b84572590608f7fb9c6db082512009630835faf6fdcb236f78e404c67"
// synthesis attribute INIT_38 of bigblock12 is "256'h2f590b4765b9de35e38e070940000820e95e950990d11d36fdba721155d0913a"
// synthesis attribute INIT_39 of bigblock12 is "256'hde4d92ae569bdb4f434fb73354cc735825a642d739f7d12ea366c7cd41be9611"
// synthesis attribute INIT_3A of bigblock12 is "256'h0dc2c7cb3b3144e704a8a00f47dcd6836d855e5b02e9d125998aa8a3cb676117"
// synthesis attribute INIT_3B of bigblock12 is "256'hff80ffffffff5039ab5c610537f284422da396ffd2f995ac4d29a5cef942afeb"
// synthesis attribute INIT_3C of bigblock12 is "256'h3a4538e6877c7f63a9af4bb02bf7f6a36ee4948103d22807b6b3fa986e461014"
// synthesis attribute INIT_3D of bigblock12 is "256'h6079ee3bba09ae7afc290b6c573d63540fcbee8ac12c5cb9946a490492c07fb8"
// synthesis attribute INIT_3E of bigblock12 is "256'hfb511d516e1ed9a5f6fff76be9e4b6c2e521dfceedfe78aaee998a18ecc455d4"
// synthesis attribute INIT_3F of bigblock12 is "256'hff807274fffb475d8770bc2a95d30a9f4cef41e7ba99b62edab616119dbbcbea"
// synthesis attribute INIT_00 of bigblock13 is "256'h597f0d98e8648ded608c2cbc6f26cd093a0c15027b771fa33e98c92b4fdb0367"
// synthesis attribute INIT_01 of bigblock13 is "256'ha8e87d1c6fc93a72b662a3471d83eec5dad28e360000801089cc1bf4dd65cb31"
// synthesis attribute INIT_02 of bigblock13 is "256'hb2b836bd62b938d934f60fd4200d5889000104005315689335bdfc52685d1d6d"
// synthesis attribute INIT_03 of bigblock13 is "256'hd65ebbae6696f417060e4ba89e7aa05dfd6b467bf4ed91c42fccbcb3d2abc89e"
// synthesis attribute INIT_04 of bigblock13 is "256'h2c10c2ce25efed17cdead72ce38657573377cd530f3c5c885608375bda1b8acc"
// synthesis attribute INIT_05 of bigblock13 is "256'ha25609162ea6e2a6e97e530d4fbf653ce6b5a6b3f30d051852e5ad95e6f952c4"
// synthesis attribute INIT_06 of bigblock13 is "256'h0580e6c01ea022342555d4f2135affff807ff800e32a558f922858cb7f7e8c83"
// synthesis attribute INIT_07 of bigblock13 is "256'hef4ac79e634acf1e27bb6db16f73854f402f27e24e66acd6cc0d400000538490"
// synthesis attribute INIT_08 of bigblock13 is "256'hac8c8a962b88df3239604ae6e41cd8a2dbe7980abf4af066290e99585a85d18b"
// synthesis attribute INIT_09 of bigblock13 is "256'h31ec49db0371ff807074fffbdee50a37aae33dac96d476d1ecb58368d8204743"
// synthesis attribute INIT_0A of bigblock13 is "256'h9f0ad7d4cd3ba3d89c38a8148b6d0087187e6ce635092e0c0d237b6723633bf8"
// synthesis attribute INIT_0B of bigblock13 is "256'h229938f9c0f53a077d1922a9d4e2a4c969533d027171b62cb7bb946d2896cd70"
// synthesis attribute INIT_0C of bigblock13 is "256'h0cc16f19aee68ca7e3a84da9aa0bab98db0074b62f659a601f992a147eb36c88"
// synthesis attribute INIT_0D of bigblock13 is "256'h83eb9541e5f388f8730e5ef590d2936e6c943b2134236f9e31fd6e6c91d1f0fb"
// synthesis attribute INIT_0E of bigblock13 is "256'h9025a526734e2c18641874cdce67b93d732f486d501627387b9450765824d4e6"
// synthesis attribute INIT_0F of bigblock13 is "256'he0ba4dc9fff9a2e6b70ef143a6ec69ccc91b833505c65440fab9fa30ee30a193"
// synthesis attribute INIT_10 of bigblock13 is "256'hc560680f428d092756884c32161a13691c91ef69a857fd0dd23be73cdf7de8b1"
// synthesis attribute INIT_11 of bigblock13 is "256'hfafd6c08393e95d2db2f9d8f2019f59f5fbee5af756d44b0d590d1839aa1a109"
// synthesis attribute INIT_12 of bigblock13 is "256'heb49b410292048177c9896aac967a7b7a8ef771fa796bdb8f2586e5d5b5f2b36"
// synthesis attribute INIT_13 of bigblock13 is "256'h9900a0fb7a10ec34dcd11551800474fffb7230ff2902c5da8e4d61474d9dbca9"
// synthesis attribute INIT_14 of bigblock13 is "256'h0011efa8ffbc1568ee3781614acc095850a36e5c9d12b728458c25734c11c608"
// synthesis attribute INIT_15 of bigblock13 is "256'h6c4adaaeb31c1c69eca392ea36efb425766e9df750c60c33aec3b4dfe391504a"
// synthesis attribute INIT_16 of bigblock13 is "256'he660675976791173d57448060149244063bd1800cde21f7028641a9d7c32900a"
// synthesis attribute INIT_17 of bigblock13 is "256'he337b9bd17efee58d5407bbc682f3b9d0ed36b029d8e403e292a16c9e5244d1d"
// synthesis attribute INIT_18 of bigblock13 is "256'hd497af967b9f0e0da351d4e8b6e1ac167581b35f231dac2e2745a6fd7d7d1d87"
// synthesis attribute INIT_19 of bigblock13 is "256'h3efb39b10c339c52f73debfad8a48c01798ef80807128b3002cb8c646d6bf2b6"
// synthesis attribute INIT_1A of bigblock13 is "256'h030e62b048009e9ba2360e7ea39952c43b68792a760ee120595fb994deb8fa9d"
// synthesis attribute INIT_1B of bigblock13 is "256'h08db42e6648639a9240b546c4bccd61795d7d74a6c9439c55d2232f2538a6134"
// synthesis attribute INIT_1C of bigblock13 is "256'h3e6bc42466d23f5d31f0ca08c55916a2ee3901158e03efbbe273a5d67627e5ab"
// synthesis attribute INIT_1D of bigblock13 is "256'h0d794c512804cd00049b682ee81bde690241000374fdfb7293ffc59bbfd9a789"
// synthesis attribute INIT_1E of bigblock13 is "256'h34ff00215ff4e9fb36739a7d167a7835681a57ef51ea548eef34bd1375608618"
// synthesis attribute INIT_1F of bigblock13 is "256'hc72d8b6a89b78f89ec9af1a9d5a1f8f2e15b968cb2ce45c70f71410cb3a2fffb"
// synthesis attribute INIT_20 of bigblock13 is "256'h494c7824b4f6faf5c97c62294a1f5df9ec14ded5969bb170200e046892dd036f"
// synthesis attribute INIT_21 of bigblock13 is "256'h166c582bddc25bcccc4a8907ddd2719378afec447f8f31134f7fdfa03033ac5d"
// synthesis attribute INIT_22 of bigblock13 is "256'he130bd0f87ca7508100336ebb79461dda0caf43d92ea54c2746a7d48d0974671"
// synthesis attribute INIT_23 of bigblock13 is "256'h2ce85ff97013bf88e2fd2c8746af41e93aaff63a321ffc18eed22c2a6478850d"
// synthesis attribute INIT_24 of bigblock13 is "256'h739542370321089a1a7a538c1828a92801021b8dbf5e25fb79e21fa554e7a8ec"
// synthesis attribute INIT_25 of bigblock13 is "256'h06d8dc28aa7b9c7111a248c34b3ef8601b57d95ba507c6cac5cb7db0490aaf22"
// synthesis attribute INIT_26 of bigblock13 is "256'h9a5f2330dbe01ba09f2a3d0f6e72880d7743d4ee3454b3ab0eeb0c87fed5a9e8"
// synthesis attribute INIT_27 of bigblock13 is "256'h9f92122044bd05734c4123a6992c649bc825861d5cd11e49000374f8fb72bfff"
// synthesis attribute INIT_28 of bigblock13 is "256'h794707af45ac0d2d2afa70f79d0e6d5914db24260000f765d40e09ff24166e64"
// synthesis attribute INIT_29 of bigblock13 is "256'hd78f20e684e0010027033f792809edf43cbe8beca9c972d894325d6bed9a0849"
// synthesis attribute INIT_2A of bigblock13 is "256'h78e508ce5ce22ee644ee1350bd6bd55afde46e8e012f45c30e52d5ab9fae170f"
// synthesis attribute INIT_2B of bigblock13 is "256'hdcdff9a447dfea609e931d54123a5028e18ec7b9d5b103fa55ca6d797cee2a61"
// synthesis attribute INIT_2C of bigblock13 is "256'hc8806732783ea5755edbc6db91241fd0a7398f26e1fdfff1bfd3b7f2b92f467e"
// synthesis attribute INIT_2D of bigblock13 is "256'h30600165cb163fd4276ed1c271a39bbb182e6ecda8981ac498544ac21ec8bd75"
// synthesis attribute INIT_2E of bigblock13 is "256'h9af8d0b255a983baa8f4e485b596cbe7960c8c64692a96dc18b1816f12905a50"
// synthesis attribute INIT_2F of bigblock13 is "256'h71b3b250b231c6b71e01ee44019d56f974e1cbe8d659aac22d50a1bbc1c6c5ae"
// synthesis attribute INIT_30 of bigblock13 is "256'h74f9fb705fff0c855f3920657ff449ddef738edf34811a96f6ddf46adce095af"
// synthesis attribute INIT_31 of bigblock13 is "256'h71d2141c6da8b3124b40433de96d0b08055c6619449b18258f445b3126418003"
// synthesis attribute INIT_32 of bigblock13 is "256'h9fdff73ba0e6c7fc8645aa5d59abb0513fab71b41ccc6b1e88db2700ef2e4da9"
// synthesis attribute INIT_33 of bigblock13 is "256'h6520659d94484280e916b142248c3693000a009006cbaad98b12ffe841fd23d4"
// synthesis attribute INIT_34 of bigblock13 is "256'h91947650d0ce3238a6747ccf92929ca4ebcd019cc40ec39895195e4ea736678b"
// synthesis attribute INIT_35 of bigblock13 is "256'hfffffdbf1dbfbffdfc865fcd14d2b7f383576e60de716223703a4d74c716607e"
// synthesis attribute INIT_36 of bigblock13 is "256'h46510010df04b875f4a6824ce10f1a3044bc956b0e3616d20000facaa97ffa9c"
// synthesis attribute INIT_37 of bigblock13 is "256'h1303436104561b8e20000120daca0202fe3e4de41b4037be43855c06045fbf04"
// synthesis attribute INIT_38 of bigblock13 is "256'h2a3ecc4cdc971b55ccab4ea1068ffdd40411de498d2d90c35d136996a864b96c"
// synthesis attribute INIT_39 of bigblock13 is "256'ha47b6f7f8991fe4d61f7faa0a9127edeac73f970dd7b6d6aa06bea69bf3de7ff"
// synthesis attribute INIT_3A of bigblock13 is "256'hd1eb41da02d2fc807274fffb36bd2b8d00294640e200e7f99732fd1f3f96ffe5"
// synthesis attribute INIT_3B of bigblock13 is "256'h0c4509e52c947c09adf04c6213ed609ca5546ac7f1257c4b24ad9b5730443d40"
// synthesis attribute INIT_3C of bigblock13 is "256'h0faf66ecfd871cf94083ba0340a865438161ab6e5465e428cd39bcf4ce9a7f45"
// synthesis attribute INIT_3D of bigblock13 is "256'h9e4cd9ca914b190f2d15e2f34ee2a3650947300217065ccdc9ac8aae9faf7c92"
// synthesis attribute INIT_3E of bigblock13 is "256'haf4f19cddd8fbc0ac4267273b5357fe6422d8dc08cff1c01a432e717d714c1d3"
// synthesis attribute INIT_3F of bigblock13 is "256'he77fffd1fd5b86ffbffeab1adfbf14743fd5f38f03f34d0b38a34be9781e9efe"
// synthesis attribute INIT_00 of bigblock14 is "256'hf0a230e09753876637605281ded6cc93e35d7256a0333e301568fceb8e76ee5a"
// synthesis attribute INIT_01 of bigblock14 is "256'h364a280096ad4000e65108c13e1051fe8a37e800b870678f1330b50560262a5c"
// synthesis attribute INIT_02 of bigblock14 is "256'h80ae8b150ade681f075470e49e88bc29449fd897a78622724a7387b6bcc31d59"
// synthesis attribute INIT_03 of bigblock14 is "256'hcddeb1e4a7d09be64ae00d684f1e0dbdd21a85e09d158fa911b172a3d7f9248d"
// synthesis attribute INIT_04 of bigblock14 is "256'hbb6a2e0454a0692f5f5b02d1ff007274fffbf63ac6fffffc51d99fe9a9ea9ee7"
// synthesis attribute INIT_05 of bigblock14 is "256'h36d480607a205815e1474269cdff3ed0b4b492ed40ee2cfa6da6e907c20a204a"
// synthesis attribute INIT_06 of bigblock14 is "256'h7430ef9c5895a02ac6c0135599f710673eb55e1aad0d5b0b9855933dcac16e35"
// synthesis attribute INIT_07 of bigblock14 is "256'h0fdd8bd915c2cb0f070f5586e660623a0a0d000022e0da01250de07433fc1bf6"
// synthesis attribute INIT_08 of bigblock14 is "256'h99fb750d393554b0dee8fcfb877e173022376bf6be84057bae8386bcfdeea45c"
// synthesis attribute INIT_09 of bigblock14 is "256'hff855367576a955f322916cd84ce67eb1e7ad105650748793485b88863a77b01"
// synthesis attribute INIT_0A of bigblock14 is "256'h68fc6d12dc74dd3b6db5349c00075be09945be99d5fe9bfa41ddff90e3fe9fff"
// synthesis attribute INIT_0B of bigblock14 is "256'hcd68502ab32600100502500150107c80797745df96b646102f1bb7a458dd02ae"
// synthesis attribute INIT_0C of bigblock14 is "256'hbbaa01dc0823bc3eeed988b29f4fe05aa449d498fa2adadf1975a439c76f6a45"
// synthesis attribute INIT_0D of bigblock14 is "256'hfeef3c5491be3d110694cf28c543d32d3596781ac424abff9bd2495be7d1cf72"
// synthesis attribute INIT_0E of bigblock14 is "256'he55b6e4b18ab9b8a2f643b7269895e5c02effc807274fffb8e90bebf8269754e"
// synthesis attribute INIT_0F of bigblock14 is "256'h6a2038db892d5562c9151010ffe6fe8d20bfffa73708288192ee60bab1527144"
// synthesis attribute INIT_10 of bigblock14 is "256'h866c1048800219173b1caabf471f6c2294de0e76353148976670d764e56abce0"
// synthesis attribute INIT_11 of bigblock14 is "256'h70f1fd9b0264c6e60ea2c1f46e1fd569f098eaf8f354e4338e313a7a402edc72"
// synthesis attribute INIT_12 of bigblock14 is "256'h3840a5246c8297efd7fa6a25fae0df3370c3529a074e5c09bb95997b156b1f86"
// synthesis attribute INIT_13 of bigblock14 is "256'hf77770f0e887f735814773aa32ff100c4d6528e61e7a180ae050b596d68b9c6a"
// synthesis attribute INIT_14 of bigblock14 is "256'h189b1dcd9b6fd62bc8b204adb6940371fffefffffffffffffd3ff9f709181a16"
// synthesis attribute INIT_15 of bigblock14 is "256'h4f93a995a8546d32002210004da6f9a4abff7ace31c94d00dda5f6930f7ca368"
// synthesis attribute INIT_16 of bigblock14 is "256'h8d356840d946864cb501f51b71bb6349e5d6263cd66945961706233b85c60c4a"
// synthesis attribute INIT_17 of bigblock14 is "256'h7a7f30be738d0e6b6b631e0b250ad0cb119fa83a5abfbed21d3ba904e990172e"
// synthesis attribute INIT_18 of bigblock14 is "256'ha07cacf16ce74d5b900c1988db6a23422dd8398b5fdb033bfa007074fffbcfb7"
// synthesis attribute INIT_19 of bigblock14 is "256'h720402da895130beaa550756ffea1c2f8f1cb072f4fe3fa7fda5adc98c910aed"
// synthesis attribute INIT_1A of bigblock14 is "256'h1448765daf6ca9060fe321710400370bab2907a337fa07eab61ebfad695c1500"
// synthesis attribute INIT_1B of bigblock14 is "256'hfd5352812455cc10dc356833ec98d08fb45411839c96aab9c2b440702c75d3ba"
// synthesis attribute INIT_1C of bigblock14 is "256'hf3145dd2d257ce8820f4fa8e83ac15de80b1f456b3b7e9cc03a7203f3410bca6"
// synthesis attribute INIT_1D of bigblock14 is "256'h9c8d0080fffcfffffffffb45f395e9bbd47f9fffdda4d9ffa55ce8750f520772"
// synthesis attribute INIT_1E of bigblock14 is "256'hf7aef33e77f08be4c60bd9d97514559ea984ca981928868d46cb705cbcbea550"
// synthesis attribute INIT_1F of bigblock14 is "256'hc50b67ac88fb3fb4ddaf1bd1f9fefd651d7333d1f37c73c5968e064f800074ca"
// synthesis attribute INIT_20 of bigblock14 is "256'h883652c16b6797db5deac0856c94dd0cdeec306ba54ae363295b6cd72df911e6"
// synthesis attribute INIT_21 of bigblock14 is "256'h74fefb729fffe5ffe7fffff1b06363a896ea92ece50caf3b1d59b92055ec32b6"
// synthesis attribute INIT_22 of bigblock14 is "256'h9157c32decc8840a54c067ad07660b25e942332502db88248d2f5989af498003"
// synthesis attribute INIT_23 of bigblock14 is "256'hb45ac4b6b3c69ddf0693dcf20d8c844aaea2216cd7156e382a02a7d02cada819"
// synthesis attribute INIT_24 of bigblock14 is "256'hd501b37f415c48fe65f276b312d800cc010000024610179c0485ef6a194eb644"
// synthesis attribute INIT_25 of bigblock14 is "256'hebfa39ea96bc52d4aae587af1937de48b24209165bc2cd2bc5e8aae22505a186"
// synthesis attribute INIT_26 of bigblock14 is "256'he64f10d34387d356764c0f4d5e5d2b21edbb5d1de928791e6989d2d79a0d37ac"
// synthesis attribute INIT_27 of bigblock14 is "256'h40b9ce205101c6db400dffc0ffffffff68ffd55d926afd9f7d4fd87765ff5082"
// synthesis attribute INIT_28 of bigblock14 is "256'h01348000265c6e75f96dd7af01f25025bf38bc8f30256d631725f63e9793461f"
// synthesis attribute INIT_29 of bigblock14 is "256'h7d672d01f672242665cb53a7a78d4f4a1338c44f5434b56832980223b92715c3"
// synthesis attribute INIT_2A of bigblock14 is "256'h648a5daa6a1ca40235a25a7a8bdec886e9a0200779cf3d3a89cc6e22d4ec4220"
// synthesis attribute INIT_2B of bigblock14 is "256'h58914e49800374fffb727ffff975757fea327a3d455bae6253eb0cbbba172ba8"
// synthesis attribute INIT_2C of bigblock14 is "256'hf8d3f3d677ff60ffc7956c4c948b514047b125620c11e9501731a2db5026eb6c"
// synthesis attribute INIT_2D of bigblock14 is "256'h3fb0767cad106a4a564f6a50d816951748dc233c244eb1750815db4b01b8ff8f"
// synthesis attribute INIT_2E of bigblock14 is "256'hcd3276c068d5265f6b0cfbac8b315713b97e0edb1e650007010402f6d43da5c5"
// synthesis attribute INIT_2F of bigblock14 is "256'h09d56b97cebc5cca14753910b082f6568fabf614fff44a9845c6d905b9a99e74"
// synthesis attribute INIT_30 of bigblock14 is "256'hf8f177ffaed4c7bfe8c44f57b9c4808b230ad4933d8a817aae079d93bf034cd0"
// synthesis attribute INIT_31 of bigblock14 is "256'hbef98d50b8dbffe0ffffffffffffffffffffffffffff88fff437f943f2f69fa7"
// synthesis attribute INIT_32 of bigblock14 is "256'h0099b1006232db5cf0af19e2fc58ee9c2cadc9e3e2920b355d89d5872829cb39"
// synthesis attribute INIT_33 of bigblock14 is "256'h59bc35a96272d20a85dbc6cfa957262104572bb44e0dee4baf215b4c29f6af52"
// synthesis attribute INIT_34 of bigblock14 is "256'hec59c0349cd95eab0c8bfd2887dfbe7842262284ff40775321688845bfaa60ec"
// synthesis attribute INIT_35 of bigblock14 is "256'h62dba027ed1658c94a41800374fffb72ffff336f5ffe480eade54bf9bc7a1e77"
// synthesis attribute INIT_36 of bigblock14 is "256'h512a0724f52cdfabf52ce7ff084297a26c4c900bb4c047ad3f620c2deb381725"
// synthesis attribute INIT_37 of bigblock14 is "256'h0c00088267f6c762927ca38269bce9fd4a32c8ca5837bd4f708ceda3a2e3ae8d"
// synthesis attribute INIT_38 of bigblock14 is "256'h381dc7d028cdbc6780a41f55f2e1a2186f5da8d1934bcf68e84d399001640021"
// synthesis attribute INIT_39 of bigblock14 is "256'h9b26b031411f51d2caa713421715fcb32e5d5b62f085771c16d5f28bf4caea48"
// synthesis attribute INIT_3A of bigblock14 is "256'hc8a23ffb157f1d9b7b94f0d55ef11a11ad77b410c4a06a70a10aa9468ed5ae57"
// synthesis attribute INIT_3B of bigblock14 is "256'h025003c8162d048426960b72fffeffffffff4fff1bde6f35847db668b2e79953"
// synthesis attribute INIT_3C of bigblock14 is "256'h4c210c0b0d4c0110004150518aa00bf9e8bb161cb480b721cdf4ad4cb83186b0"
// synthesis attribute INIT_3D of bigblock14 is "256'h908eef25888d8506dbff80108624f7ac12e17d6042d21f557fef465a795cab64"
// synthesis attribute INIT_3E of bigblock14 is "256'hf8488ee3b221302437b4bda3cfada1e41b8dfd9c7eea071fe9274c04bdde7c45"
// synthesis attribute INIT_3F of bigblock14 is "256'h0b69aba0133022db30230c3dd8b39b41800374fffb70f9ff4d7f5fd06cffdffd"
// synthesis attribute INIT_00 of bigblock15 is "256'h93a46b0fcae302212c889f12db6cbfecfe9d087fc7966c4c8d0b54c0a7a53f62"
// synthesis attribute INIT_01 of bigblock15 is "256'h00120040000028021d3277fc3d22cb7e9a0544744c1c15de56ca185ac48581b4"
// synthesis attribute INIT_02 of bigblock15 is "256'h524512b9931f23c1db736623de33b13156ac161ca4874fce263d904676b366ea"
// synthesis attribute INIT_03 of bigblock15 is "256'h24b2dd4806265426fd4ac7b53d3b87fef6b77bb5bb8658f1cd500622d6a97aff"
// synthesis attribute INIT_04 of bigblock15 is "256'h153beff4ba9da2611afe576a1413daafcff5f409aa7040b91b9c21e8d1a8a772"
// synthesis attribute INIT_05 of bigblock15 is "256'h3eab43544c8d824360c2eb82963971b6001380002008da0674e5bf20e3c17ff1"
// synthesis attribute INIT_06 of bigblock15 is "256'h8c8387f284f4028a2000020122001a20acb1fe667b4e6ebed1bb79396f419513"
// synthesis attribute INIT_07 of bigblock15 is "256'h2360e9d5a4c250e07dea6168abc859d493ed8fda2f3474f9ae1191b2f341ae0e"
// synthesis attribute INIT_08 of bigblock15 is "256'hb2147bffffbc3dd8503f32a0278f1d7dc048513e2f2e0e1b8226a11d195c44ad"
// synthesis attribute INIT_09 of bigblock15 is "256'h48852c5566e6b9754a0b1927db33220246a8c1ed425903a7ff807274fffbfffa"
// synthesis attribute INIT_0A of bigblock15 is "256'h3767e51a240064b18d6226e300086068e65829aca5bfa90f17fcad90dc918b6c"
// synthesis attribute INIT_0B of bigblock15 is "256'h859120361161200800000140129b97fc5268b51b80b3770745cfc2a3e523595d"
// synthesis attribute INIT_0C of bigblock15 is "256'h348c9028e738c1aa1e8810ba94232d4ec9426603ed296d71304406d90c04a21b"
// synthesis attribute INIT_0D of bigblock15 is "256'hfe8c1afefacc56319ed6090065697776f93bf2a0464bbc78806b12506bcfe3e8"
// synthesis attribute INIT_0E of bigblock15 is "256'h7d03e8a5dccb5126767d2736851bd6966b1ab91bff01fe8fafeae9fcd0bf7fff"
// synthesis attribute INIT_0F of bigblock15 is "256'h4f60c1e126ee5cee52d1cb5a1646d6579083098fa1920400c1c2bd9c7e8520ed"
// synthesis attribute INIT_10 of bigblock15 is "256'h3abd47996ecd80372885ec72a51dc7e762e4bf1a4fb883fc06cbfd3e43baec66"
// synthesis attribute INIT_11 of bigblock15 is "256'hb6e7a16a91d03d278a37465ec9655aaa7a19789c4354c53c4bfac8adc9048589"
// synthesis attribute INIT_12 of bigblock15 is "256'h7274fffb51bc5fcca7c5b15bd937d94f389f3d03ec99262991f3dd5fda26ef90"
// synthesis attribute INIT_13 of bigblock15 is "256'h2d51e8938aec408dacf467a76505200b2569db3d26c23f18e1ed4f59038eff80"
// synthesis attribute INIT_14 of bigblock15 is "256'h9bb442df3ae8c4fec711d41a5e6130ebb06da5119c6d0104608437dd14ea1a0d"
// synthesis attribute INIT_15 of bigblock15 is "256'h37b1240b186ff69b14146296990e4001006bda002a9408caa9b42756fe69e885"
// synthesis attribute INIT_16 of bigblock15 is "256'hfa782d67077e1b6bb6aeb74b0bb6824c7cd8161511e4ef5b52c5cf92155c662c"
// synthesis attribute INIT_17 of bigblock15 is "256'h26a01b2609ad93ddc4519b62fe36bde52635e4c2aea5d5c7888bae316a60bb6d"
// synthesis attribute INIT_18 of bigblock15 is "256'h0044bfe8db524f754e830281db852c191fee817d79414ffbe81ef7d57de97d77"
// synthesis attribute INIT_19 of bigblock15 is "256'h2810a6608dbcad8f0392e236a64afd60aa83660124963673d4a113216db510e4"
// synthesis attribute INIT_1A of bigblock15 is "256'h8446262396c14e780e01d8e903f70bd49b2ba51589a182c742dc70ca44860000"
// synthesis attribute INIT_1B of bigblock15 is "256'h4d155ae33dbc51b98a209af82108d0045c3ad365defe66c8cc7698e010fae58a"
// synthesis attribute INIT_1C of bigblock15 is "256'h415a02b8ff007274fffb7bdf5119b7b875498224ab9f46f8ec7c090ff7df5545"
// synthesis attribute INIT_1D of bigblock15 is "256'hadeafd20c6f7a4481c910b6de095317368a6893d620f24c7db431c825480612f"
// synthesis attribute INIT_1E of bigblock15 is "256'h08c499a89c5ba5de66525a61717c942db6fba1056d60b8dc0168f24aa63d889a"
// synthesis attribute INIT_1F of bigblock15 is "256'h5487fe4053280e1749e347bfe55e98d95b59be3b00060042829065e0f5aa2db1"
// synthesis attribute INIT_20 of bigblock15 is "256'h4fde7acd2aab1ec14ddabaeb6c98c7bde28b2641bfb2341fe339722fb24add69"
// synthesis attribute INIT_21 of bigblock15 is "256'hc673346edddf1f12937bb30abf69363327b9149abc2ada50a30716755642f968"
// synthesis attribute INIT_22 of bigblock15 is "256'hffffffffffffffffbfff70a15653d402e24bfad22f0cbf8fafe6246b65f5ed9e"
// synthesis attribute INIT_23 of bigblock15 is "256'haf7d8044b9d2128c6ae7da8211b4b5b38e8c0c0cc8323a596d50b7240140ffff"
// synthesis attribute INIT_24 of bigblock15 is "256'h7529e6db21319bb56b87dd1afaa523a573e9a8a60c2501590000b134e718037e"
// synthesis attribute INIT_25 of bigblock15 is "256'he528c1175a038f272196a039155144106cfdc48a8407274e4e7085bceb1bb650"
// synthesis attribute INIT_26 of bigblock15 is "256'h20021798c9eb485a0383ff807074fffba16f77ff7e554efda163557f43935385"
// synthesis attribute INIT_27 of bigblock15 is "256'h225b4d0083879a9fbfd2ca7e89695cc50aede088ac536ae4953d644c24c7ab5a"
// synthesis attribute INIT_28 of bigblock15 is "256'h63851da06c803f8a93aa62ce4bd7188c58f5eb48547a95eaf28fbb78aa1791b6"
// synthesis attribute INIT_29 of bigblock15 is "256'h417e801054dda0df5f96c28726bc442f91012b236a5796078aab001009800000"
// synthesis attribute INIT_2A of bigblock15 is "256'hea464d518edd07c37df5b94e9b6331013c3f42eb06239f426a385f51623b9ade"
// synthesis attribute INIT_2B of bigblock15 is "256'hfffffffffffffffffffffffffffffeaf4ff4f6fef5375229ddd93f92f7744224"
// synthesis attribute INIT_2C of bigblock15 is "256'haa96161360ea0183ec39b4b0402a4264b60f8f1199c883eab582dc6d0124fffc"
// synthesis attribute INIT_2D of bigblock15 is "256'h5ed166fcda7301fdc955589d34a60abdc9be9a41257b176e5080e4a696eef292"
// synthesis attribute INIT_2E of bigblock15 is "256'h567fa4c74f46060e5d9ff3511e5e1ef7fee204189db540eabdd95840d6289bca"
// synthesis attribute INIT_2F of bigblock15 is "256'h14c3a86cd256e664fb6ad4c86de03e9c79db129c542abd689ca15fe9e0f5d404"
// synthesis attribute INIT_30 of bigblock15 is "256'h0a752d1e373182dbf823ec5a59b1d048800374fefb72d1ff13999c1b3ab3f655"
// synthesis attribute INIT_31 of bigblock15 is "256'ha13d36da006ed00159cfe9fff2a0a67fe4a498afc4896cdc8b8bf64067a00566"
// synthesis attribute INIT_32 of bigblock15 is "256'h9590836dc0114ac65ddd7e508c6e60c079c23ac2d52190aa38a5cab4f4bec81e"
// synthesis attribute INIT_33 of bigblock15 is "256'h95ca193365b6fcc3c913979a1fcdd05ea9118863a0add473448d49aa54e5bfb4"
// synthesis attribute INIT_34 of bigblock15 is "256'h9f2aeb18afcc0fe97beacca9eaa823668e604f99c6f8d4f213871ad315e506ff"
// synthesis attribute INIT_35 of bigblock15 is "256'hfffffffffffffaff57d77f93f949abef8a40edfe17ce37adac2373be8dd71500"
// synthesis attribute INIT_36 of bigblock15 is "256'h568f20a4d10c06ad181b8d225925d212a5511c6dff81ffffffffffffffffffff"
// synthesis attribute INIT_37 of bigblock15 is "256'hb8ea3e50c52e1ca43f49c67a025c5d0f190af1102c4212de69d3ed04d97fd726"
// synthesis attribute INIT_38 of bigblock15 is "256'h565f63154191619187d2d7bbb60cb9bf1166f01a8a562533894121444b36b236"
// synthesis attribute INIT_39 of bigblock15 is "256'h6fd5532b79bb273e4c9b52018a6f7d6e254b30d982d94d56d94e9032d3600e59"
// synthesis attribute INIT_3A of bigblock15 is "256'h55a027ad3d660dbd2b80372442db30258b6dd9c90e32800374fffb7275ffe91c"
// synthesis attribute INIT_3B of bigblock15 is "256'hee013103220a1a484a0806c3b6d6037157d2abedd9f6ff2889dfc31decdc848a"
// synthesis attribute INIT_3C of bigblock15 is "256'h84999cf8a8e3327f00110400060ada22e974dde886a1c5e14eefe423b6b60135"
// synthesis attribute INIT_3D of bigblock15 is "256'h9a11ddc962dbafb08b7cf52f780835be87efd30b7456fdc1a1d4699e90ec2da7"
// synthesis attribute INIT_3E of bigblock15 is "256'h77fff5775dfb7634bbb7d475d28054bcbfa64074bfe0f9c4c100a00115aa205d"
// synthesis attribute INIT_3F of bigblock15 is "256'h0803d31a69f229137fd0fe00ffffffffffff5fff7dce0f3557fa5bbdff92f96f"
// synthesis attribute INIT_00 of bigblock16 is "256'h10cf755148658694117ef1c1f1d025a5fbf80b8ee41a53e438223ca3600b9383"
// synthesis attribute INIT_01 of bigblock16 is "256'h6bb4ac914bce1589eb2452f9c3e96817b31e2b87796b32ca000096400be5c463"
// synthesis attribute INIT_02 of bigblock16 is "256'h3f7e2e20efd9a80d488cf67646f000d56b2cfc864da97634b45b2ef85d8477d7"
// synthesis attribute INIT_03 of bigblock16 is "256'hfb72f5ff6b7ffff58a96fffdff98696f8dda793201f5c8c4cae52fec3c4a9340"
// synthesis attribute INIT_04 of bigblock16 is "256'h94946c4c908bad0007b107624b7de8901331e2bb9024ed56d8898948800374ff"
// synthesis attribute INIT_05 of bigblock16 is "256'hf3969be5b3068435b9adc6310b8da8cb02bcb8d4028de64aefe32979fd91f8ff"
// synthesis attribute INIT_06 of bigblock16 is "256'h4abc2f72051b918ddd190dad818d04d482006a204d1eda666a5d3fbe10ad958e"
// synthesis attribute INIT_07 of bigblock16 is "256'h5893b9341c2c8ae80f847520f2f01a1e57318b5a7625bdc9a9e31111ab859976"
// synthesis attribute INIT_08 of bigblock16 is "256'hc015e930a467fa680ec617903129feebfe9089c110aaa9dd8506371d23761227"
// synthesis attribute INIT_09 of bigblock16 is "256'he040ffffffff970ededf60694c207f4d60c2fa7e0ab3d7e8239bac2327ad674d"
// synthesis attribute INIT_0A of bigblock16 is "256'heae142dfcdf9187cc1786a5a781e264b0ceebf503253c5c12bb50a7a8da986e4"
// synthesis attribute INIT_0B of bigblock16 is "256'h25dade95b48dff46aa43555b26a0040bf06bb948333f585300000012c0006800"
// synthesis attribute INIT_0C of bigblock16 is "256'h88d2fac2a6128769a330c5e350dd423ed8c886229bb21c2b6125658e9a0e58fc"
// synthesis attribute INIT_0D of bigblock16 is "256'h0748800374fffb700fff4aeebfc5fff24656effffb20be6b2a1f1a54a9a6fe63"
// synthesis attribute INIT_0E of bigblock16 is "256'h2afd320ea8ac66346c8c8c8bf84867a477640c216768222504bb1030e23e5919"
// synthesis attribute INIT_0F of bigblock16 is "256'h17a74a34066bfb416a347c1977ec25af17ad0bb89141db6b0938c0000ac07dd1"
// synthesis attribute INIT_10 of bigblock16 is "256'hd6f1636515662d9410eec2e991c0986b6eabdc61400101009047f68cd776a7e6"
// synthesis attribute INIT_11 of bigblock16 is "256'h1ea6870af3f3c630da25ddd9a8a422913c3bfbb065be9e52dd7a5c33bb5a0b54"
// synthesis attribute INIT_12 of bigblock16 is "256'h3eafeff7c4ffeafc3357eaf7f65d09e6f40c694f17458625bab82b286af30fe5"
// synthesis attribute INIT_13 of bigblock16 is "256'h582c50dfcc5e541b4af99d17620c4094aa7a71c6045bbfa8c3a25bba15ea2852"
// synthesis attribute INIT_14 of bigblock16 is "256'h2dd1d68b76614db4a54209b6ca6257d2d33c01510010e4000794b3e75ab002d7"
// synthesis attribute INIT_15 of bigblock16 is "256'h605574172e129563f8ec0490ffb53d856844c0b12b6080105b03a5774fdc6ad8"
// synthesis attribute INIT_16 of bigblock16 is "256'h113db0e130507c4e8a2ca89604812a85240cbda206ac700a496f9486962322e7"
// synthesis attribute INIT_17 of bigblock16 is "256'h22a23d58b1ed4fd9038bff807274fffb3a0b401470f04aa13c8134f512950c7e"
// synthesis attribute INIT_18 of bigblock16 is "256'hf1f77bf547eadee11e2a173d2da0e8c40b6c008f3d5267a6c9050e0b1928db37"
// synthesis attribute INIT_19 of bigblock16 is "256'hd1304ae1d8d12541072859cc1b6d51b90007d7001bb6633d64b9f14f69cdbdc5"
// synthesis attribute INIT_1A of bigblock16 is "256'h90e5b468bf6d5a726247e79ecb8719162babaa5e615c32962461000e01406ac3"
// synthesis attribute INIT_1B of bigblock16 is "256'hdad37144acf559660f5b6369d7ca0f5a2dd46914d6ad218be5da66b3d05910a8"
// synthesis attribute INIT_1C of bigblock16 is "256'h331194cf555433b143c31ec0aab44bb90b3ba0c36d010a5cf65cb366bca55743"
// synthesis attribute INIT_1D of bigblock16 is "256'hc080ffffffffcbafc495fc64b8ff455df5aa558f67f76be91baf319ad6b03d6c"
// synthesis attribute INIT_1E of bigblock16 is "256'h47db7da528fe01c82040000235b25ad91fb8b7c620384513882a6a88c91b0371"
// synthesis attribute INIT_1F of bigblock16 is "256'hf5f559284923d3b449bcb9d9b9f7b881dcfaaf6f2cf724069102d201ae633623"
// synthesis attribute INIT_20 of bigblock16 is "256'hd913851d75c2ce973553d2c77f0247d39afa2431f0c0aa3f55f6784b115a35eb"
// synthesis attribute INIT_21 of bigblock16 is "256'h66102507db571ee26d28c9e9485a0311ff807274fffb4398fca2277ab9d5ccf3"
// synthesis attribute INIT_22 of bigblock16 is "256'h896e102092c727d6fe9122efa7f4ea3bcdef0c89683305adc853b1096b47295b"
// synthesis attribute INIT_23 of bigblock16 is "256'h040b0022cf00054447fd67e520446da9c8d6387ec8363d735c441ad8566646da"
// synthesis attribute INIT_24 of bigblock16 is "256'h2b656b313923eca49e6b666c8d458d8a6bc8ab8b1f38ae3bd4f82379e366d533"
// synthesis attribute INIT_25 of bigblock16 is "256'h4cd61d1f01a1cccbfdbff532f9f1de8b9e2f19f31eabfc1fd2fdf2beaef52178"
// synthesis attribute INIT_26 of bigblock16 is "256'h8148bd0417b95d2e44b75b6f5e3e9422a0b832f79bd356570c37a054bbbd8fd4"
// synthesis attribute INIT_27 of bigblock16 is "256'h97d936b51b8efff0ffffffffffffffff751fa6347523916a5be1812d4ffa58f9"
// synthesis attribute INIT_28 of bigblock16 is "256'h32cc10000c95990bd07b67484c9eaec81afdd8fab0ffd68f5dfa060c25a838a4"
// synthesis attribute INIT_29 of bigblock16 is "256'he8af5f2422679426ac36a1529a3e63ab7f1c8216a9e7c96243138fe5b51985b1"
// synthesis attribute INIT_2A of bigblock16 is "256'h7e99d555784084afb229913d3c2681ff54f1058b4415c733d53164c9625004fe"
// synthesis attribute INIT_2B of bigblock16 is "256'hacb56b279d5b044c0cc64b5a15c14628b1ec565a03e2ff007274fffbb5baa43f"
// synthesis attribute INIT_2C of bigblock16 is "256'h0e18641513e0e0c7da446e36c5404fffca7fdbffff43226b1ce85c838b6d6078"
// synthesis attribute INIT_2D of bigblock16 is "256'he954c45b31b006b0480064008502391f3f5c038d4768fe0c9aaaa19717ae3751"
// synthesis attribute INIT_2E of bigblock16 is "256'hd0665676a18030ea719d286406a4eead766850dbad29302ce880f4d33c8f20d2"
// synthesis attribute INIT_2F of bigblock16 is "256'hde25ad5f04930d8cec846e6130beae83f1d77ea318fe01599878c603bac91d30"
// synthesis attribute INIT_30 of bigblock16 is "256'hfff0ffffffffffffffffffffffff27fffc89a6fffffefffefffdfe3e917f7ebf"
// synthesis attribute INIT_31 of bigblock16 is "256'hf9fd8eb99578abab752327d17f626d238759e45a4311406a4ddbd30a8e460403"
// synthesis attribute INIT_32 of bigblock16 is "256'h376a3c37e9a5503b8d64411b49d32f199f8e18f3a60bc000202582753d7a1105"
// synthesis attribute INIT_33 of bigblock16 is "256'h2f3983e589253e3cce15217990e9fb479b5cc182726215180cd4ec64c7b196da"
// synthesis attribute INIT_34 of bigblock16 is "256'hfffbf975fdff37a8df537313bd73f39487a43d9bb736dc8a9a58a1fc4eba8b0e"
// synthesis attribute INIT_35 of bigblock16 is "256'h8c650b6c4087b14d64476923900a31e7db232282471811ec48d903f4ff807274"
// synthesis attribute INIT_36 of bigblock16 is "256'h6b55a539d8a1ac40b6fc839b54c838479458db502e38acb8f9efff397f5b9cf8"
// synthesis attribute INIT_37 of bigblock16 is "256'hd33c1891ba413fec4f068cee4dab3aef100043ae7e755163667e184bc551ab2b"
// synthesis attribute INIT_38 of bigblock16 is "256'hffb29350062e4552ba8d895430a9bf4a23b591b3f2c40dbd51fc32eb8de3234a"
// synthesis attribute INIT_39 of bigblock16 is "256'hfd5b03359a84c39f325ce8202d518e84b6c702a1705946fd53c7133f84006032"
// synthesis attribute INIT_3A of bigblock16 is "256'hd2426e36ffc1ffffffffffffffffffff883f9577eefd5677fb7ee367fcef538e"
// synthesis attribute INIT_3B of bigblock16 is "256'h672078f90c94ed84a2a6b990add1d9b78ee98ceaf0eb496984d958f8e3b34885"
// synthesis attribute INIT_3C of bigblock16 is "256'h4d158e40c29357f00521088b60352f5382d8dee654d7c4a2775a7ba211c80000"
// synthesis attribute INIT_3D of bigblock16 is "256'h0a5a994373b2abb1d075b29811943a2563851b33e452690e3fbbc62006c99a7a"
// synthesis attribute INIT_3E of bigblock16 is "256'h0354ff807074fffbfacda5d7cc13b75a24bfe9296b3950b210252c89e9c4a5e5"
// synthesis attribute INIT_3F of bigblock16 is "256'h297f15bbae084cc78b6cc091adb462c7e905900b31ebdb1726e25482b1f85e58"
// synthesis attribute INIT_00 of bigblock17 is "256'h821dabb43b401e404d0bbb34946eb87c4fa28a37b4c1dc6d4800f133b2b3ddf5"
// synthesis attribute INIT_01 of bigblock17 is "256'hee0d2ace78c1a00b93ae8d281a7de72ba6b9c4ce000401401d127f349b5dddd4"
// synthesis attribute INIT_02 of bigblock17 is "256'h44ffa1342fd6b62932fd362d3fa2473d8f69970747ece88be9fc629db4c3a3fd"
// synthesis attribute INIT_03 of bigblock17 is "256'h6df96ead301b61f7236e199dfa4aecaab4176e66b22fa648a21e8930ce32935d"
// synthesis attribute INIT_04 of bigblock17 is "256'h609726a8abc45b7f57d647beddda07fdffe3ffffffffd227f46c2797feba6baf"
// synthesis attribute INIT_05 of bigblock17 is "256'h5120802087cad02675ffffb18925303807f21683d419d080f13fe7e7d6383153"
// synthesis attribute INIT_06 of bigblock17 is "256'h579a598ab45cbd48498e4df8a35e4937e224512f5caa26b929195f15d36d010c"
// synthesis attribute INIT_07 of bigblock17 is "256'h547245bf417e8e82074141f2f116cd3bc1b7c7a27443f97c85100524a426269d"
// synthesis attribute INIT_08 of bigblock17 is "256'h2023095558936a48800374fffb72b5ff91710d129c187f66ddfbf29f6ffffffd"
// synthesis attribute INIT_09 of bigblock17 is "256'h441b636c441d5ed845549018c2b56c4c838bacc06c3105620c85e7581325c2db"
// synthesis attribute INIT_0A of bigblock17 is "256'hc953f4111c2fecb798f1113c42f93231280817101f543062e6a9371c90424b33"
// synthesis attribute INIT_0B of bigblock17 is "256'h20033118d8d55a901086f11da3c0603be58453a40dd4960a42a0001100008f22"
// synthesis attribute INIT_0C of bigblock17 is "256'hed283be49217cf4878f826b638040688de3d4ce58812090bb4643f7a19a8c595"
// synthesis attribute INIT_0D of bigblock17 is "256'hffffffffffff8a7f83e0dbf839ff09fba7d195d3f6bf1a5b2faafacb2b064f28"
// synthesis attribute INIT_0E of bigblock17 is "256'h10eddab603f2315bcfabd3431d3ac9140ea91d1a2b2a6b14da626eb80000ffff"
// synthesis attribute INIT_0F of bigblock17 is "256'hdd0dce4e0902365d5e4b02364c51b0592081e0528af279e16829000608049472"
// synthesis attribute INIT_10 of bigblock17 is "256'h17ff4ad7f59b217f3446c373ab7bee24888c275ac35d4c63e2f9e98576d52070"
// synthesis attribute INIT_11 of bigblock17 is "256'h47203630463d59f5005cd289cdffe26cbdfc5b0819fd6f26c6d8ef76418ae964"
// synthesis attribute INIT_12 of bigblock17 is "256'h6868323cc49b582ce96bd9b13b4f800374fffb7270ff65ea675450b45e9963df"
// synthesis attribute INIT_13 of bigblock17 is "256'hb6ba1c919e826ce8c41e177aa0895953a1d1911decccc3934cc0e7b103660a21"
// synthesis attribute INIT_14 of bigblock17 is "256'h00260480a694e4e8c2c2bdb50720e21584158ed53d16f35651a622508d452369"
// synthesis attribute INIT_15 of bigblock17 is "256'hc6cfaee6692b11e15b621573d72292a4c3b34799783a4520326975cb00183400"
// synthesis attribute INIT_16 of bigblock17 is "256'hefb8de1d2a9efa443affbc3814a77bf8b62e1cff7efec5e5d8aeee19af5fd0f3"
// synthesis attribute INIT_17 of bigblock17 is "256'hef52d21fdeca826c84afa9f4732397b913b455be1144bfc9f4f7049276d41ee8"
// synthesis attribute INIT_18 of bigblock17 is "256'h83172f173083839c5548c6db520d0002fffeffffffffffff2fffc74a7328bf50"
// synthesis attribute INIT_19 of bigblock17 is "256'hbdd921483007e2cbf70d1ed1a52c12d4031d00000bb07f08fc9c18689341b916"
// synthesis attribute INIT_1A of bigblock17 is "256'hac1cab5584c71d1fbbedcdae856e561fe9bba9c55d72b3b50033291a77a2c5db"
// synthesis attribute INIT_1B of bigblock17 is "256'hf18435c05cc16c33688af9d4575e94d403055d4aeba35acf6f5b0396f6b5deb9"
// synthesis attribute INIT_1C of bigblock17 is "256'hc63d23640ead654a272542db2020e953d919ff41800274fffb72e6ffdecc71e6"
// synthesis attribute INIT_1D of bigblock17 is "256'h6dac16e4280026007a5e95b195fab9e48232fa75b10cc842919d6c8c820b53a0"
// synthesis attribute INIT_1E of bigblock17 is "256'h55a55816350c000280800910a7f2dbf4031ff906c7a47aeac1b00c9dce93daa8"
// synthesis attribute INIT_1F of bigblock17 is "256'hf678520b095d818f133ddef59ca113d9a69f37cacdd3fdc2bb6037409c57f2e4"
// synthesis attribute INIT_20 of bigblock17 is "256'h654ec0a9543499a9714872ae235ad5747fe514d41be3d9c152596fdbf34bad9a"
// synthesis attribute INIT_21 of bigblock17 is "256'hffff390fe2c24f44fc58e21711d99fbb96057e884cba9a3cdf7a476e8f85574b"
// synthesis attribute INIT_22 of bigblock17 is "256'h424274e0f8451a2f73aaa4b5b5996042091e0761f2e76244358cdc8e2102fffc"
// synthesis attribute INIT_23 of bigblock17 is "256'hdfc4d4ababf4bbb66e7a7b32a762ba28cdf844e4c8dbd482ca78011b800008a2"
// synthesis attribute INIT_24 of bigblock17 is "256'hedf101a4783447f587a49dbb5e34a0d47b73b7a66fe62e0b8d48195f99717c61"
// synthesis attribute INIT_25 of bigblock17 is "256'h1dfffd058593a884adabceeedc75d152c6ef3c049ff896b5cc8bc504ae58e5f4"
// synthesis attribute INIT_26 of bigblock17 is "256'h2de8700b5e60e620216e0d5d48387a0c41fbd81a2f445be99f41800374fffb70"
// synthesis attribute INIT_27 of bigblock17 is "256'h65c6ec588533d6abd97236d60b8e38200d003d70cde8aa7ffffde51d403f648d"
// synthesis attribute INIT_28 of bigblock17 is "256'hc4315acfca3331dc24b800c4000000002f4ae1035bb3fedd97a85412f1a8953e"
// synthesis attribute INIT_29 of bigblock17 is "256'hf08d83cc8986b80d54db409f97f0495f40a2935d3151924313b484aad85dc1b6"
// synthesis attribute INIT_2A of bigblock17 is "256'h808ef46589893fc7dceac048c7c03914ccf928723e2a667f7fccd84999d1ce60"
// synthesis attribute INIT_2B of bigblock17 is "256'h8cd5ad17d8eaeb54db540dc6c100ffffffffffff4bff961edc2d2dfee5fff137"
// synthesis attribute INIT_2C of bigblock17 is "256'h595ce86885589b2e135902480000f8b98c83ba70e81af941b32dc08f2706ba4c"
// synthesis attribute INIT_2D of bigblock17 is "256'hcdf36a7218648e4a471faa36bcb7d8ff690f7b8072efa55158d5414b26704f09"
// synthesis attribute INIT_2E of bigblock17 is "256'h3d3ae9250c1065514d09603137c6174eee29aa5434fff39cc3bf8fe5ec6e3fed"
// synthesis attribute INIT_2F of bigblock17 is "256'h0366ff807274fffb9caf0249deaa8d314cd30e09d7131ace66aa0e97361b715e"
// synthesis attribute INIT_30 of bigblock17 is "256'hb13da69ba52068b18b6de87facf86ae76173900d2162db571e622f98b9e740da"
// synthesis attribute INIT_31 of bigblock17 is "256'ha6a33654055d99215c052b69b3d68914f6ad07ff588084f0a63ad15e4807d7fd"
// synthesis attribute INIT_32 of bigblock17 is "256'he6f3b1eb66429a242ac2b272ccf1b36d4347400244809200036c898a0c32e250"
// synthesis attribute INIT_33 of bigblock17 is "256'h7f7288b3ec4b73c05f2f2431030aeba440b4d008f46b24d6dcc2f68c11a8ffe5"
// synthesis attribute INIT_34 of bigblock17 is "256'hfffb6fd62ff92fff434be8ff5c97fce1e8d4084ed96ec673a4cf01a9c789effe"
// synthesis attribute INIT_35 of bigblock17 is "256'hbfb5da0c544003ecc6a55a8dfff0ffffffffffffffffffffffffffff9fff387c"
// synthesis attribute INIT_36 of bigblock17 is "256'h498d0bb27ad9895d001b01008834413839bff12335f9a681ae04e2468eeba5b8"
// synthesis attribute INIT_37 of bigblock17 is "256'h2d3ea533c7459699666fdbd763e25c532d436ad56ebb0b4c95a2313b83751a8b"
// synthesis attribute INIT_38 of bigblock17 is "256'h4eb891e2ba163833193ccd3e3527e09beb858d8fe8b9759f24a5763a5a2ae1fd"
// synthesis attribute INIT_39 of bigblock17 is "256'h3c60d1eb3259031aff807274fffb3f9c5169b6df4576b73004f406a1f040e2ff"
// synthesis attribute INIT_3A of bigblock17 is "256'h08bc7f9482cc99ec9f141d10d8f3092c2079b4fe6647893b664e2d05bb372042"
// synthesis attribute INIT_3B of bigblock17 is "256'h7b9dd0bda2907b721923739d42eeff100381ca91942e6a1eb71c06015828bb91"
// synthesis attribute INIT_3C of bigblock17 is "256'h0544daa1d4d0e043513d40e518d6f29149d9c9f71a9339a999e15bdba0007e0c"
// synthesis attribute INIT_3D of bigblock17 is "256'h91fc2ba1d490727a3bdc8ba56395298926ea46b7ba89c4d496da585865de0d43"
// synthesis attribute INIT_3E of bigblock17 is "256'hfbaf015ba7d5661fe0c9ccf16d6a68217734316f35954313638f61f03f1fb596"
// synthesis attribute INIT_3F of bigblock17 is "256'hffffffffffffffffffffffffffffffffffff2cbfef956fde3383f442d33fa1a3"
// synthesis attribute INIT_00 of bigblock18 is "256'hcbe14c4e38916500d24a62d951789f54c6bb92468d1ca81ce391fc16ffffffff"
// synthesis attribute INIT_01 of bigblock18 is "256'h097116d64d528dcd6cc98810f8099f17b7b8f438c24e52920fd30011c0805484"
// synthesis attribute INIT_02 of bigblock18 is "256'hc310a459c7ae210ffd647ee7834157902bd0b756e2f03010af36c26922c559b6"
// synthesis attribute INIT_03 of bigblock18 is "256'h1988db3320425530b9e940d90354ff807274fffb37ffd3e6047f7fc33ce66d75"
// synthesis attribute INIT_04 of bigblock18 is "256'h371b0041fb05efeb2fffdfffffa0e2fe2921cc640aec2078acfe66c7a921360d"
// synthesis attribute INIT_05 of bigblock18 is "256'h124000400c1536640602e7bdd412d4948ec99902e2210629f8d44f3806a16945"
// synthesis attribute INIT_06 of bigblock18 is "256'hcb10708af5f0f475e7118ed25895b96e06ba9924873afd1eae82c649babcbcc6"
// synthesis attribute INIT_07 of bigblock18 is "256'h44eb3ebd512ff50703ebc6a4052a38128ccbdb2690ca904e1401d53011c54f94"
// synthesis attribute INIT_08 of bigblock18 is "256'h8b7ffe9f340befeafee72dfbfa935d7f1125eaf4e21fd4899cef82d4c0c497f9"
// synthesis attribute INIT_09 of bigblock18 is "256'habb9c1de3fb9b21c0f9eeb815b9a8a68deb422360ddf49eb291bff02ffffffff"
// synthesis attribute INIT_0A of bigblock18 is "256'h42a95791e67c42d1dafc0d42ae5b8e7200558000a5408f8384df3ac27d3ac9a4"
// synthesis attribute INIT_0B of bigblock18 is "256'h442c4c50a8c8269e53ea386cdea9e1099e9cf8b78460044c4a7f620fa3175939"
// synthesis attribute INIT_0C of bigblock18 is "256'ha95f54c05f7f24c8eb30e56f3c9980e799696b406de60114a449b34f63328d17"
// synthesis attribute INIT_0D of bigblock18 is "256'h6667b1771c0a192adb331dc255c889ed4f59040eff807074fffb9b7b44d2f529"
// synthesis attribute INIT_0E of bigblock18 is "256'h93b6c905a2fcb4ff8cf16d4449233d007f5ae9c3ff3d9560dc960b2c4080a855"
// synthesis attribute INIT_0F of bigblock18 is "256'h16f57bad6ca410010a002f0c2c9089db3b19815fa5168736bba3a2e31aabfd3e"
// synthesis attribute INIT_10 of bigblock18 is "256'h4ccb7dd579ab6378d41a25f9e2ac6b59ae79e78adbda8d89d57c7c4839c86161"
// synthesis attribute INIT_11 of bigblock18 is "256'h02423427a8c732ebebb57412a38037eee8e66aace166dc2e6b3cbadff75a0951"
// synthesis attribute INIT_12 of bigblock18 is "256'h62ef90a252f506ad08189944ac43b86ca1a49f7294cd32bd82a6f48a2eb7e81b"
// synthesis attribute INIT_13 of bigblock18 is "256'h7c93b3699d1959be02512b43001383c1fec000ff95b0fbe7bfc757b5c554fa1e"
// synthesis attribute INIT_14 of bigblock18 is "256'h8ad4b70c2403c41d9717382d000208005124402ad50495745e9ab832e7a0a07b"
// synthesis attribute INIT_15 of bigblock18 is "256'haa105222839956eaf1eea951040961db08be8833e15edf97f364b26e538dba22"
// synthesis attribute INIT_16 of bigblock18 is "256'hfffffe5329f5799773fb5c62279a34ca166607c0f22dd0601f19f0342c539369"
// synthesis attribute INIT_17 of bigblock18 is "256'h6c0c928bacc007b125610c45caa0033c42db1026e86d58294849800374fffb72"
// synthesis attribute INIT_18 of bigblock18 is "256'h1fbb3a53319eebb1c0c0f088e5b87c67a6d7838db200f4aeff5b4dfa90eaf4a9"
// synthesis attribute INIT_19 of bigblock18 is "256'he1f76c0cd608d5e4a95a02e821c01f5e8b12f88480d3e64746f4c126d512a246"
// synthesis attribute INIT_1A of bigblock18 is "256'h8d4b2e543ba12945a80efd617c293e03f0f740e56461be35f8e1ddef8fcfc0f0"
// synthesis attribute INIT_1B of bigblock18 is "256'h88556d519bf73116de4443ae496928c1b480ce2b5c7c14ad80acf571f1b205b4"
// synthesis attribute INIT_1C of bigblock18 is "256'h91b416dc1d0400c06a7ff50cb69319be189a57639faaf21337a70256d4e29f37"
// synthesis attribute INIT_1D of bigblock18 is "256'h3200894901429c0a228da62662fabba1799484d685a204218be43ac5460e9108"
// synthesis attribute INIT_1E of bigblock18 is "256'hdead85bbb528ba4b8129484a604423b2011293a56507a901602101d32a810000"
// synthesis attribute INIT_1F of bigblock18 is "256'h7193eba1ba665ab54609331e7b966aab14faaf1b93c967ab68d8f1e04752b814"
// synthesis attribute INIT_20 of bigblock18 is "256'h800374fffb72b6ffafd0ed0fdd2910d0b8142579d7dd01128b8f22241b7dfa6a"
// synthesis attribute INIT_21 of bigblock18 is "256'hdf4f084dc6ae6c9c960b5200263d23650af9e7282619a2dbb823ed2e5941a957"
// synthesis attribute INIT_22 of bigblock18 is "256'hc085246891c9715bc3006b8271999894d72ea3c1eb3c91738a19e34f623fe262"
// synthesis attribute INIT_23 of bigblock18 is "256'h7b04eb8490d2dc37a4914419000001197d950620943dc8f55d61b06248c36afb"
// synthesis attribute INIT_24 of bigblock18 is "256'h6ad3adb33292069510b52ed4b7ab8f79f168a248c56097fb3a85ec4a44f568ce"
// synthesis attribute INIT_25 of bigblock18 is "256'hecd95f945469d61b9c9e7e908dd8802b874253785c38f9af8d37fbb8b311f875"
// synthesis attribute INIT_26 of bigblock18 is "256'ha1c3963fe392584858c0d8fdb10bc2a16ac66919f63a013c1602ffaef54ad4d0"
// synthesis attribute INIT_27 of bigblock18 is "256'hbabcbe3b049f8f658da017c53c936850b91b0371c451ff255fca287cebca075f"
// synthesis attribute INIT_28 of bigblock18 is "256'hdd58419a4bdea736531d76af63331786a8cb407022e307af020000100005174a"
// synthesis attribute INIT_29 of bigblock18 is "256'h799075d4113900916ba55f72110e903a5ec252c8c4156a81973d7b10d7a8080f"
// synthesis attribute INIT_2A of bigblock18 is "256'h8f545b494050800374fffb72dbff1fb733fa59d3546d9df4ffc8d4ac0797a34b"
// synthesis attribute INIT_2B of bigblock18 is "256'hca00efffd494ff7b89cd66182da86306136044bd256d0edd272a6d0d62dba824"
// synthesis attribute INIT_2C of bigblock18 is "256'hef5e3404cc8eda52267b0d5e1674a8d3c85fe3241c460fd7da36723680002804"
// synthesis attribute INIT_2D of bigblock18 is "256'h22a992ef2baf3484eecacd5d29146821939455dbdb4c0002000102032023a5b5"
// synthesis attribute INIT_2E of bigblock18 is "256'h458aaea491f7b3a49da2904734ede5ada8001577d807ebf1fd30a07c1ec42791"
// synthesis attribute INIT_2F of bigblock18 is "256'h7ffef51fd49fada95fef46a60de559a290d062244c9069e5bf9589c75e1fbea4"
// synthesis attribute INIT_30 of bigblock18 is "256'hbe0e746793d6ef083f655e5f694cc8db0001c180ec0fcf76f4bf59e83fd5a77d"
// synthesis attribute INIT_31 of bigblock18 is "256'h85168515f2393656800500000d0088f0ef40405af44c098f8b12a75be979e5a6"
// synthesis attribute INIT_32 of bigblock18 is "256'hd6187765c3cfa70bdfaa304a34839438e9b315de4dce1312bcfe287114754ad5"
// synthesis attribute INIT_33 of bigblock18 is "256'h673ca45743207903a8358f9eb6208aa0fd2760f06a3e7060088a8fe53abedcf7"
// synthesis attribute INIT_34 of bigblock18 is "256'h4a30416b7818ef3cda41d24e800374fcfb709bffb31d9a7335538cdf7a09b13b"
// synthesis attribute INIT_35 of bigblock18 is "256'h86ebbeae22247fcc4bd975f38cbf28f2f4896d34978bed0087a43b694b152360"
// synthesis attribute INIT_36 of bigblock18 is "256'h5b457476c5ff27d5e971f3d75228644e62d111a6779d6db400dc000000c07509"
// synthesis attribute INIT_37 of bigblock18 is "256'h73cb15505e77b06a1ce3a19c946df91b109c200080002150c2b390af10f8de7f"
// synthesis attribute INIT_38 of bigblock18 is "256'h7e092140b258899b4541c599de0b0d4719b81539d6162e04cc7db71487991a33"
// synthesis attribute INIT_39 of bigblock18 is "256'hf388cda1a2fe4b6e6aba2b331f9cacd59be84e0bda9a57c96299773de2513dde"
// synthesis attribute INIT_3A of bigblock18 is "256'hdb4ce695cf5dd7d2a43cb44d9dcd6d91352300007850d951ea3bfc8ff51fbfea"
// synthesis attribute INIT_3B of bigblock18 is "256'hd856e751941c1caaeacb0034000020020e040507376b3d54103d08601d3ef72f"
// synthesis attribute INIT_3C of bigblock18 is "256'h3e2b5dc3966ebfacfa87ff04a7fa0492421af9e9b0a159a4910c729d5049c903"
// synthesis attribute INIT_3D of bigblock18 is "256'hdd7d02ffd3e59a8651113d561fa076451c0658ac5a6fbc7c5848c4d1ebb35cf4"
// synthesis attribute INIT_3E of bigblock18 is "256'h658c913d4a4d3d25bb2a25426bf049eb4ed9033afe807274fffb1dfe7f54f55e"
// synthesis attribute INIT_3F of bigblock18 is "256'h8e6a0f93236d0037480083bcbdf9e8df97ffd7ffbf959561b4f40aec8098314d"
// synthesis attribute INIT_00 of bigblock19 is "256'h14c00a005b80c511064f8aad632b83831d41cf1de1c842b9c7f4768198b98098"
// synthesis attribute INIT_01 of bigblock19 is "256'h54cbf3995460954799e58e974a7e450d823382507f228d47953eb91f504825b8"
// synthesis attribute INIT_02 of bigblock19 is "256'hdb70b2bf82a3f10accfffcc41b557245e88d7ab7e158d9880c40510e8aad3d69"
// synthesis attribute INIT_03 of bigblock19 is "256'hff82f6cd51001be8fa0e1febf303cabfea046fdbe94ecb3ea8510f95980b373a"
// synthesis attribute INIT_04 of bigblock19 is "256'h00a5ea8bb9d5925d9650a81a89dc2350d4da8913c24d1a0c72470000f8004715"
// synthesis attribute INIT_05 of bigblock19 is "256'h35b6fb0524417076f4582a61aa75f94d5150a00000000d61d351f1c7319837cd"
// synthesis attribute INIT_06 of bigblock19 is "256'h1a8f1160bb0bb1565ef19964478a75b64d114ce72dcaa04a4a0de3ca5f4918f1"
// synthesis attribute INIT_07 of bigblock19 is "256'h477fd3f3479bde8c15fe2aa2156da723416190067245bcc744b1c0700dd57d64"
// synthesis attribute INIT_08 of bigblock19 is "256'h8aecc0959c5a65875977580c3d65db2a24426d3061eb47d90315fa007274fffb"
// synthesis attribute INIT_09 of bigblock19 is "256'h7078422a398894ee08d88a5d8ad98a878db6005bbd41c7e789b02ceeac39a8f4"
// synthesis attribute INIT_0A of bigblock19 is "256'h7d352dc92922477c13370731004011d3588232db586312cf403213332d533398"
// synthesis attribute INIT_0B of bigblock19 is "256'hb6e7bf5f75ebb9484c8ddebfe378af8c313da0dacf75d9eb415238b9e59c8653"
// synthesis attribute INIT_0C of bigblock19 is "256'h8c13db40d39eca9450efb9204425c8973e6bd40da1011fe6f376a9f58783b82a"
// synthesis attribute INIT_0D of bigblock19 is "256'h0009004006fea22af5b3e82b22fa7a9cb6bb083461c1ca379d473f10b7a039ab"
// synthesis attribute INIT_0E of bigblock19 is "256'h2c89d819a8aff7f6767915c25dce3ba179b760aeb7babe8ebab43d9b4f9ac6e3"
// synthesis attribute INIT_0F of bigblock19 is "256'h34d053859add6588b3a01ea216d70f6ca88e1838664ca26996246866452a2025"
// synthesis attribute INIT_10 of bigblock19 is "256'h528c3332b655e4179c0dc1fad34c9a1f186380e275ac164a518b51a182897658"
// synthesis attribute INIT_11 of bigblock19 is "256'hfd807274fffbf51c3bd73d2efb20aabb3624bc4eadfd0a1347c5cb4fbe240540"
// synthesis attribute INIT_12 of bigblock19 is "256'h171ab4204cf40b6c8096c1526327e5051e0b3d2ddb1a26e215c0b30b4858033c"
// synthesis attribute INIT_13 of bigblock19 is "256'hf8947ad454d3b02d48f224a524be03eb248d04a99902f28225bfffa32a67bfaf"
// synthesis attribute INIT_14 of bigblock19 is "256'h68dd5a58dbd72544ada611da995a0521010120c000102631dff4e5376fef6802"
// synthesis attribute INIT_15 of bigblock19 is "256'hc7e1de5fde37aafbec290821da11e66d6ac2f8b70b397015eeb96a23e9064bd1"
// synthesis attribute INIT_16 of bigblock19 is "256'hcea7d6e66abfeb346fff9945d6da27a9db2365f028323e7316a4ac9e5bbf6e8f"
// synthesis attribute INIT_17 of bigblock19 is "256'hb8a1b6604aba3525e2b40549e4894136ff00ffff7fff37f47674fa676dfaffce"
// synthesis attribute INIT_18 of bigblock19 is "256'ha15661d8fad374a6304700a1a560f0197da0956d86ae0da20e9eb9e469262a37"
// synthesis attribute INIT_19 of bigblock19 is "256'hd2b34ae75cf798bbfaaa1248dd49ad6f44b186a2606946f574a5a8c99e36df2d"
// synthesis attribute INIT_1A of bigblock19 is "256'h7e8e9d310d169a3c122616c45ebf301d0809d4a5cfddd6276f5fba443e84e7b5"
// synthesis attribute INIT_1B of bigblock19 is "256'h29eb48d9034fff007074fffb3185b7e6731f3a15fa1a1ea9c24aff9a11673a07"
// synthesis attribute INIT_1C of bigblock19 is "256'hf0d74d2f3476ff33ac109cb10b6ca87cb4f364a40975820d31a8db2a22e23f18"
// synthesis attribute INIT_1D of bigblock19 is "256'he31a6a82b5c5c620bb82b42ff85a35184acb90261b8f8b9d050d49a682dc66a5"
// synthesis attribute INIT_1E of bigblock19 is "256'h4015b3d2671266b6465696f611c31067562b197e6b2b2347300000004075c2c1"
// synthesis attribute INIT_1F of bigblock19 is "256'hbd8c112e0860120b972ae2de10d3f413a8b04a97208bb76f81b280b83440be0e"
// synthesis attribute INIT_20 of bigblock19 is "256'h7fcf8d9eee4073b1c7f37a87fec0fb9f97a8cd2107ee70a79d4ca802e506a36b"
// synthesis attribute INIT_21 of bigblock19 is "256'hd2ca78c42c68349003515f4ed673655d83e8efbf5ff5ed74afffb5dd93f3eadc"
// synthesis attribute INIT_22 of bigblock19 is "256'he490012200000900f248175ffc6a835c540094de5cca2370af26a12e98e5c875"
// synthesis attribute INIT_23 of bigblock19 is "256'h552b0e4c33cc3096fb552752d1a1648cbf2701342537a95ea344fb98ff9bb492"
// synthesis attribute INIT_24 of bigblock19 is "256'hc1ea1e086d93b1958ae2bd5d10e2117eef0f39d2f56e06376a0fe2dcec6c1bd3"
// synthesis attribute INIT_25 of bigblock19 is "256'h172502db40248f6cd8d1284f800374fffb72b2ff210b1bb017cfbc49ca7442c7"
// synthesis attribute INIT_26 of bigblock19 is "256'h69a72fb669101240217a7f9fed104076b7966c4c878bf360263c3f620d65ac4c"
// synthesis attribute INIT_27 of bigblock19 is "256'h55424315b1de3f578f13b243fbff2ffa0a3653c6db9c463e8342356275dcfb50"
// synthesis attribute INIT_28 of bigblock19 is "256'hfffbe9ffffffbff7ffbeebffe99db4599b66ffd5dbffffacf9ffcebfad965994"
// synthesis attribute INIT_29 of bigblock19 is "256'h6b11511433156c5275d92e4f9ae0652842f4226effff3fffa060c0aaebac6fff"
// synthesis attribute INIT_2A of bigblock19 is "256'h5106f3d5fcd44ad41bad7054556ce39a9f79a48899d34b0d89b40e523a5d624d"
// synthesis attribute INIT_2B of bigblock19 is "256'h8ad5403de4fc8fe397bc903942086067e595133197a300006a00109132753db7"
// synthesis attribute INIT_2C of bigblock19 is "256'hd4f17311695dd5558e813284464b324c753856462445c974f05ca07cacc89559"
// synthesis attribute INIT_2D of bigblock19 is "256'h8b0a4a08132464c34b55c759a46430279290bc9cb09717669470a3541a6c4531"
// synthesis attribute INIT_2E of bigblock19 is "256'ha06ba71f939f06bd4429d8495229fcbc2d7bf979bc37fe64eeffc52809e85c55"
// synthesis attribute INIT_2F of bigblock19 is "256'h855e154d2c00f3a642ca08233d6057c58f50800374fffb72d4ffffff0fffe8fc"
// synthesis attribute INIT_30 of bigblock19 is "256'hdd4c4a051aade3fd113143d4f8f79afefbf514bc00c61ef02bcbfe0f80005997"
// synthesis attribute INIT_31 of bigblock19 is "256'h6a6e6ce63c5b4f47000b83004ac9ab73c6240dbec6234b45b73459ace74ec601"
// synthesis attribute INIT_32 of bigblock19 is "256'h7dde82c804c4165a0710863a238dc58966b59f238a3adba0fd9de4dc6152ff6b"
// synthesis attribute INIT_33 of bigblock19 is "256'hab4a2f38c6eca50af0b4815b9323889279d56d194c0e72eaded18deece6268fa"
// synthesis attribute INIT_34 of bigblock19 is "256'h659b6526994a9dfbdfb643bc719c279fe4c91b71e250e9301ab5acbdf09759ab"
// synthesis attribute INIT_35 of bigblock19 is "256'h516db295d8e0ea4dd85d397aff04800fb658abe29298c69075825969ce280277"
// synthesis attribute INIT_36 of bigblock19 is "256'h225a3872e0057a486b652400ad5bb6ce4f0460e73e34de0ec437cf69e6666a9e"
// synthesis attribute INIT_37 of bigblock19 is "256'ha997d43e682ed114a101154fd623403867be53bf5bbab4bd8c4384018234faa1"
// synthesis attribute INIT_38 of bigblock19 is "256'hfa01755f516654784f8338266263503b7e6875f40b7f8b98876000d9465a283a"
// synthesis attribute INIT_39 of bigblock19 is "256'h920c0020dd8611644f8d240022c663ab002e6520d916d640000374cbfb726dff"
// synthesis attribute INIT_3A of bigblock19 is "256'ha9390964fb8eb1223ff06db74b6b5db30059dfaff3fffeb707db012c8c806c8b"
// synthesis attribute INIT_3B of bigblock19 is "256'h026b4f1624df49e8b9019eb23b3aef2047737d16674f6f87bf5dd32f0486e796"
// synthesis attribute INIT_3C of bigblock19 is "256'h182331288279034a2eed58f5632dc1ec1b5c5a1528e7a5923be9b69b3f8e8dea"
// synthesis attribute INIT_3D of bigblock19 is "256'h091e7066cd4afcd45ee8b595d824fd91973320a487325e5db2e69c6ba1fbb412"
// synthesis attribute INIT_3E of bigblock19 is "256'h4013445f0dc2b7d8236db5e7c665ab062c3b7f1b528bb4d961650fb1b9e9e48a"
// synthesis attribute INIT_3F of bigblock19 is "256'h43363cbfd1257668b6ecfb0a29fe48d634eb8f558bb469b5f2e41db1d26f08cc"
// synthesis attribute INIT_00 of bigblock1A is "256'h6ca41546271475bbe545097406c86f424d0ef1bdff91d6c3a140c1f9d9a448dc"
// synthesis attribute INIT_01 of bigblock1A is "256'h97222359d88bfe17ca42023d0dc14d09b33e991511fafbac73c87d5cb6f9ac53"
// synthesis attribute INIT_02 of bigblock1A is "256'h74b1fb70dbff91b659645c52f5001f81850bd1a7d01defa32aa6f373334c7e7f"
// synthesis attribute INIT_03 of bigblock1A is "256'h293e2199efb490086be0a618fd7d4becc390ed0ca2fb5a23281bdf69a81e0002"
// synthesis attribute INIT_04 of bigblock1A is "256'hde9b5b8dee11e7987fd438d688c3f298097724abcfd0611b1a58f7020506e181"
// synthesis attribute INIT_05 of bigblock1A is "256'h630e9471315cd1abe7dcf1d234c0046ad9e42ab302f4a759a3101eb89d146c00"
// synthesis attribute INIT_06 of bigblock1A is "256'hb83c4ac4e45de0a53181d2ebe363cc756d42b8e0956623af532edc95d5eba118"
// synthesis attribute INIT_07 of bigblock1A is "256'h101a760e6c9cc6dbfc8d9022d6444a17e8e097dac5d4286b14624a1b190becfc"
// synthesis attribute INIT_08 of bigblock1A is "256'h902935b822930c26745b88eefeeaa6558a826d995333144b70e398e0ba26bb41"
// synthesis attribute INIT_09 of bigblock1A is "256'h59271205d4424e6a7a3ac10d8b0bdb65ad56412f8ad94d90a679506702cece71"
// synthesis attribute INIT_0A of bigblock1A is "256'h02263a2802a874b186acc1f533a401493983a139c788b47045878bad7188b532"
// synthesis attribute INIT_0B of bigblock1A is "256'h7ac1d593c1e39f4db6d39c29003681091409628c4cb9a62624bd5c4f96a1f52a"
// synthesis attribute INIT_0C of bigblock1A is "256'he923535f02f1bd807274fffb4a83d615d5f2a458a07071c0b189de222285cbe6"
// synthesis attribute INIT_0D of bigblock1A is "256'h052904da952904c49518f42090ef6098047e7fa4f8ff244a04430bfd24031658"
// synthesis attribute INIT_0E of bigblock1A is "256'h64a0f0c20fc3503ebd5a185cb4ee198aa73edf8e09a9a496408bfd60f6aaa16d"
// synthesis attribute INIT_0F of bigblock1A is "256'hff19912c8e64655ddf20b6a4ffae9c589bfa8306081abe3bb782ccf82e95c5f1"
// synthesis attribute INIT_10 of bigblock1A is "256'h1fc63c266cf9a6db5d70c3da7fe3df9ded19fdad08bb4fef6fc0f8cfbbd528b3"
// synthesis attribute INIT_11 of bigblock1A is "256'hd0007126caea8ea53d84d1b7feeb723b2958f8cc489e0c851822c7eac373603d"
// synthesis attribute INIT_12 of bigblock1A is "256'h2ae303b1986159b1748816f6e3f292f54dfc8e0dac1d8bc2ace2d86cc57b2a72"
// synthesis attribute INIT_13 of bigblock1A is "256'h502918b34eb13050bba899f94679e5960bf80d6661c432e9eb5288ad314c2748"
// synthesis attribute INIT_14 of bigblock1A is "256'h87efb0a9ff85d4ff4c78a47f908628e1a28c3358ab859ae8ae43f5c4a5e50d30"
// synthesis attribute INIT_15 of bigblock1A is "256'hf28d810440e3942909a7ad8a3f461b7615d9b4ad3dfd24c7c806ea6e42733d9c"
// synthesis attribute INIT_16 of bigblock1A is "256'hdbdd244231e0e8c9185e02b9c8807274fffb560695cbb052cb6a804ec45cabcf"
// synthesis attribute INIT_17 of bigblock1A is "256'hd383d18168a348297fcf75ae64c30c9968130aef0893206f7ba67c87440b0c28"
// synthesis attribute INIT_18 of bigblock1A is "256'hb340d3cc9628110e6c7769dac8852f783eeb60fbe5cca634c36da9e4b3cf94c9"
// synthesis attribute INIT_19 of bigblock1A is "256'h11a3a860b8ed1b6d0e4748d2cb72685caf14fcb05b590513334ab825b40a9d42"
// synthesis attribute INIT_1A of bigblock1A is "256'h2926428a0b25f4124b8de47b28ab3a392604095c5332af71d058e92f674526f5"
// synthesis attribute INIT_1B of bigblock1A is "256'h5058acebe359eda99f5bb0c6ad944d442212e1b978b1a43fd9f51760a9485004"
// synthesis attribute INIT_1C of bigblock1A is "256'hb9684866f0e5fa44397beecd68cd43e92d620e21eec8648711035feb1902f505"
// synthesis attribute INIT_1D of bigblock1A is "256'hb8dbca723122c7d0cb9a85c8bb3b9ed831c4de9189c511650c72c8de291877cf"
// synthesis attribute INIT_1E of bigblock1A is "256'hdcd2770a7ea5d273a81b6cf61629be771e7c489b5fd960ab2b83466269c06da7"
// synthesis attribute INIT_1F of bigblock1A is "256'hacdf7d53c0ac726eff5e57e0d411cbe843c5c5554864fb3457ef939eb64046f5"
// synthesis attribute INIT_20 of bigblock1A is "256'hfcbd260a04c22be920e41b286989346002e7d5807274fffbe5ffb07533dcd6bf"
// synthesis attribute INIT_21 of bigblock1A is "256'h3a3468af1ded5ab906cbcb55210c0057d55292398db2b46290f1c0a1a0747da4"
// synthesis attribute INIT_22 of bigblock1A is "256'ha450fbbd7effff4b950821dd9dcb474333a752c73ab4fa7a8590936cdcb2cad4"
// synthesis attribute INIT_23 of bigblock1A is "256'hd0003fd542774987d6ac38370751288004c6b419b6d75c6d52c7189c2b447790"
// synthesis attribute INIT_24 of bigblock1A is "256'h636980c35537976eca9b19710017651c444566838743a0731d5b0125cb4d1a5f"
// synthesis attribute INIT_25 of bigblock1A is "256'h95443f4cc16f0907d6dc57613d5f45015af11c2aab790ad52ce61829b8aec3a5"
// synthesis attribute INIT_26 of bigblock1A is "256'he26b8f48fcf0c5b450df6de1ffdae1be1574faa178e785a29c7a3eaaa53f7b18"
// synthesis attribute INIT_27 of bigblock1A is "256'hdaab7b26a45a9d0053f56db4c9db43756b442b4e16eca5b62687a5a49c401678"
// synthesis attribute INIT_28 of bigblock1A is "256'h59a6282080a545248b411e1602044d8757633cbcb74fbba53b505ec570cbd1e2"
// synthesis attribute INIT_29 of bigblock1A is "256'hce701bad4f8c6255d40efa6e01d40fd209215a05a12e6b5beded01c445aaa44a"
// synthesis attribute INIT_2A of bigblock1A is "256'hc89eb0497fa7316da20c08c23bfd24a41d10e928415d02f2e1807074fffb7a11"
// synthesis attribute INIT_2B of bigblock1A is "256'haa48fbf274672acc7d9dad179cc610f99a31b6bf8e7c528e954d0a18f42490ef"
// synthesis attribute INIT_2C of bigblock1A is "256'hc2724ca846a26da636dab56f40ade41159e3469cc76c21a95a52c41698693197"
// synthesis attribute INIT_2D of bigblock1A is "256'h481e0017889808250060e8db2a7ec2ba98b5a6ef4827af7eaed4744cea16352d"
// synthesis attribute INIT_2E of bigblock1A is "256'h3c85e657f25ffe06ccb4a5e5baae48d96cf493b7355a634f7cbe16802c2b9b6e"
// synthesis attribute INIT_2F of bigblock1A is "256'hdeb65bb1395ececedbd4c9f272f9d16f916226779b43306f20ed100d6cf6ad65"
// synthesis attribute INIT_30 of bigblock1A is "256'h6fff19915e0466926b3447faeb3ba9e2ba0944b85094300530d8db9f1996e71e"
// synthesis attribute INIT_31 of bigblock1A is "256'h590f36a21763a1b1175157b11aebbcd55acc943872a6b664398b9a460b64792c"
// synthesis attribute INIT_32 of bigblock1A is "256'h0d1aee91e8f44668dd2f345831edcb62123308f1e025c90a6bcd00da09408951"
// synthesis attribute INIT_33 of bigblock1A is "256'h74e6fb72c1ffcd428bd5de8ae617cf0adaf15bd565f29e9998b68399af44c58d"
// synthesis attribute INIT_34 of bigblock1A is "256'hc187578aefa88d8d5640a324ff7d0b3ce35e0d18243c2827881de07915430003"
// synthesis attribute INIT_35 of bigblock1A is "256'h5818b3c55890ce5815bd8e38397388732648ef1a59519160ccdc7442e8fff228"
// synthesis attribute INIT_36 of bigblock1A is "256'h70e1a38ff91a266a6aa0de3a4d8aa0e087a24a1c7308bfff822a48c81d99b5aa"
// synthesis attribute INIT_37 of bigblock1A is "256'hefd6ab8d8cb11c9d514a6d53c701a9d52239c5aa800595c89e83221b2d6cf592"
// synthesis attribute INIT_38 of bigblock1A is "256'ha7159041572ac7dbd982ea555a9b5cdfc2be779df925f3d1e769c26a189999e7"
// synthesis attribute INIT_39 of bigblock1A is "256'hdf68c4fd3d62e7449deebab165f5acc8559e9321115ac3f2df4102bbcc8d3112"
// synthesis attribute INIT_3A of bigblock1A is "256'he93e8171383a8eaa50e25daeb620d36d4a98fad4bb2128c66f41c5bf7d01f636"
// synthesis attribute INIT_3B of bigblock1A is "256'h9833faaa2ac094005729b243ec48728602b8597ba324073fe445f83adf0f48f3"
// synthesis attribute INIT_3C of bigblock1A is "256'h53d41458329106aa4df9563589364799db9f67a5a0e94d4426360e01da346590"
// synthesis attribute INIT_3D of bigblock1A is "256'h5ce9263b800374edfb7219ff9de3bf2ca943b83ebeb258d3b8e730f7674f1dc0"
// synthesis attribute INIT_3E of bigblock1A is "256'hc2b649ff2da6001d308aee64858a750044acd7734c30c5389904641ba0242f34"
// synthesis attribute INIT_3F of bigblock1A is "256'h67206dcfa4db12ea482cb7199c0651587f258bb90dc9136a63495814f799d4b4"
// synthesis attribute INIT_00 of bigblock1B is "256'h2eac0881e36b371dfe891a2f9ea9940dd2b6453fb6559434de621280ad3b40e3"
// synthesis attribute INIT_01 of bigblock1B is "256'h3f238fa0229e6d3102486d0e7c246a07e691df94e6de4f8ca09cae2ff23502e4"
// synthesis attribute INIT_02 of bigblock1B is "256'h867c836c9b53caa5a24cd32854cddd900874da3db3be1a500ea4dc40e15f3be4"
// synthesis attribute INIT_03 of bigblock1B is "256'h7d07fff7382ab7afdeb3739cc8351154e868aaf2a7302d67e15d7f437a1ae556"
// synthesis attribute INIT_04 of bigblock1B is "256'h75d23702238abcf01e72616acede8c89930002ccaad37854275b48218611d818"
// synthesis attribute INIT_05 of bigblock1B is "256'he3363d4b7ecf167a1621e29b83d91ad194a3c8e0ec920b116c74d38add5ec001"
// synthesis attribute INIT_06 of bigblock1B is "256'h85e780651a040d544f7596a8b2477d92acaf940fc608f3ffc748f55306b26a1c"
// synthesis attribute INIT_07 of bigblock1B is "256'h443b90288f2ddd51334b800374f2fb7295ff071f434fa8e9aa9c28f042044b38"
// synthesis attribute INIT_08 of bigblock1B is "256'hc9a1b481cb94de764105169b91d730a5eea8958a78c0449411750bc16594aa09"
// synthesis attribute INIT_09 of bigblock1B is "256'h2f9816b51e7a87f047f6fbd9c0938cfbdcf68c098846b8322ee37fff90db0ac9"
// synthesis attribute INIT_0A of bigblock1B is "256'h16f56b79fe96cae5d6d39042455362385919005d001940012600b28a31c95a05"
// synthesis attribute INIT_0B of bigblock1B is "256'he6ad81849776a54688f67133a1ff40de17561f4cfab4735ef8908c5f75e58ab4"
// synthesis attribute INIT_0C of bigblock1B is "256'hd239d2792fcb0f2450b99e46547295b418a11b7b77d6a20dca6596703a07f998"
// synthesis attribute INIT_0D of bigblock1B is "256'h5dca11ca46992309b4aae08d05f700007f81b9bda8b1490aac2420b51f1f65f6"
// synthesis attribute INIT_0E of bigblock1B is "256'h2c2511c1a64f66d3029800ac03008d0e21f98c2dfec3d735f509d1cb18c68aa9"
// synthesis attribute INIT_0F of bigblock1B is "256'hb41a2506d7bee4c097d9217175c98fa8a89246b8d6245ec231fa53bd07a8eac1"
// synthesis attribute INIT_10 of bigblock1B is "256'hf6bbd25f8f415ea722138b5b61676b8f8167d47935e166add11d435857851628"
// synthesis attribute INIT_11 of bigblock1B is "256'h0c44a266960c043b402288155cc9f044800274f4fb7010ffc103a7560a253745"
// synthesis attribute INIT_12 of bigblock1B is "256'h988affed026bb2b4736ea98ff28e7038142c51a723166e5893901600463da573"
// synthesis attribute INIT_13 of bigblock1B is "256'hae0e477bce597f3b16fdbca5c0605a37f4400212b8d44616620ddac30684f986"
// synthesis attribute INIT_14 of bigblock1B is "256'hb3ab97c19373032890d3e549a8769596598d142bea6a8ee83d113d80502d61c0"
// synthesis attribute INIT_15 of bigblock1B is "256'h24a202a9d2e2aed86c99133ff79a6fd73d6290ecd621389f51ccc318c1d1a63e"
// synthesis attribute INIT_16 of bigblock1B is "256'h4807cddc8c568755bfddcff2877b6dad668fbeb65f7c2ec932925ec6b516f23e"
// synthesis attribute INIT_17 of bigblock1B is "256'h185e2ce72c9ba842f6b36dbf18db4229891267c05ffcefbbfd6c93df2ca6e85d"
// synthesis attribute INIT_18 of bigblock1B is "256'h0eae8f1094e2dc0005b642810d24663d4181c18cf7afa14a64a03abbd431e942"
// synthesis attribute INIT_19 of bigblock1B is "256'h12e98e336352ae4317d2bed6337db7a8904e46be7f1aa4873f97f6067959908c"
// synthesis attribute INIT_1A of bigblock1B is "256'h4cc26d5d39329b5b53212e487fcda7bfa4e0e797cb1657374309d6cc6f16272a"
// synthesis attribute INIT_1B of bigblock1B is "256'h009abd166f2570f5264c05259b7922e31e30e1e84bdb0341fb807274fffb9e5b"
// synthesis attribute INIT_1C of bigblock1B is "256'h659e36db1a67a0227009aefa96a1735bdb4cb8263557ba0ed3d02da1d8610e6d"
// synthesis attribute INIT_1D of bigblock1B is "256'h0e45258fd13f0fa9ea58ad5b042bab41b8dc1af6be13fbd43c20154710b76a0c"
// synthesis attribute INIT_1E of bigblock1B is "256'h98feabe759df7f9f5c82a238ff5c8475567b0ca81cf9e38806a8a00069281a00"
// synthesis attribute INIT_1F of bigblock1B is "256'h9cf9aa9da185b8aece2714009e33edbd168167d57f839f8e54d8b8eb65636a9f"
// synthesis attribute INIT_20 of bigblock1B is "256'h35b91841ceb7b3668bceba765cd14b5eae7b98a35cdf64bd8fc92cdaf5945fb5"
// synthesis attribute INIT_21 of bigblock1B is "256'h48b4a4cb2de048a856db506dc297f86bd7a90ad4fd905efbafdd79e76f6b089c"
// synthesis attribute INIT_22 of bigblock1B is "256'h089734939024e818ef8cd2f6a961d5bc8c76b099aae2348346cc14df0fdfa506"
// synthesis attribute INIT_23 of bigblock1B is "256'hf9f838ef7ead2a77e604ad53308ecd4708f72737ce3b9c5b5a8aec23ad2a1c37"
// synthesis attribute INIT_24 of bigblock1B is "256'h7274fffbf33f5c8854363907aa24e83a356bd58a9c1dfa155cec3481664873b7"
// synthesis attribute INIT_25 of bigblock1B is "256'ha621b432106ec0a2ac7675a4e511664b18a29bad262332fa61eb445d036afc00"
// synthesis attribute INIT_26 of bigblock1B is "256'hffe68bbfa3b8a7af98e486852ce9c677c3a8f2e250811f17a377fb0b72cbe062"
// synthesis attribute INIT_27 of bigblock1B is "256'h0195f88f85494c42f518d05a35d557e3d4c5a8cfa5a9e0f7271ff356147008d9"
// synthesis attribute INIT_28 of bigblock1B is "256'hc5674e590b21c98a87c426962c23f92f2f0b60d3b54f89234c3d001998a01292"
// synthesis attribute INIT_29 of bigblock1B is "256'h53d191dc4546f92b74f25a8fa953f356913996b9ca177f442726cffa0039dd6c"
// synthesis attribute INIT_2A of bigblock1B is "256'h4117adb3657ddbc8895a48a8e673eea4302b673b49b795a365184ec8cec886a4"
// synthesis attribute INIT_2B of bigblock1B is "256'h809c0c0c67c926b776e56baf1d460794309c3bf36db78a63ca0c2162e5fba851"
// synthesis attribute INIT_2C of bigblock1B is "256'h95d4f2a67fffe0106aceb58758fd26742029c8e0194e65243c5fccc9a935ffe0"
// synthesis attribute INIT_2D of bigblock1B is "256'hc9a0a38322b684900ab83f14d06e7acaa3d24130f16b663eb11513f92a10a794"
// synthesis attribute INIT_2E of bigblock1B is "256'h43dd039af9807274fffbd6962a24d6aa62ed4315a82dd35e84db4b437b7fadbf"
// synthesis attribute INIT_2F of bigblock1B is "256'h5303231bb58e08a1a4138eee408f147a75a6b8f72a4b04c7abaa26234caa692f"
// synthesis attribute INIT_30 of bigblock1B is "256'h71fbb6da238a451494093246e48def4d22721d4520d784eb6aca8ac98a98abf8"
// synthesis attribute INIT_31 of bigblock1B is "256'had631364a489561af074f0a171bf2048a47fe39cf5027a3674af065161e5e6b9"
// synthesis attribute INIT_32 of bigblock1B is "256'h1f4d163dade7d2711d8807d67f9775efe0573579a8a9eee48a3128cae8008d3c"
// synthesis attribute INIT_33 of bigblock1B is "256'ha33ab68d0ef2fbe39739f81d1a929ae93c6e58f16635136ce84de456d2f18d80"
// synthesis attribute INIT_34 of bigblock1B is "256'h089ca278508a458b8c7fc7393ba8f9dfea43d9ecf5aba7411def54b2e8c56cc8"
// synthesis attribute INIT_35 of bigblock1B is "256'he1218745723e70141b169be2b22a9ece82f6a6d8ac004401b7de336da0bb1198"
// synthesis attribute INIT_36 of bigblock1B is "256'hcf5b9699a8b91b3b233df1f77b48c4f64151755026a40a76112d718454467295"
// synthesis attribute INIT_37 of bigblock1B is "256'h7f915280eadaf26e4b83fe12304cd6bf41e4eda3fdd6342cdfeecab84ad6ce64"
// synthesis attribute INIT_38 of bigblock1B is "256'h2404154a692b585e0330f7007074fffb13f0f429cea1a5bcfc5ec23b820565de"
// synthesis attribute INIT_39 of bigblock1B is "256'hcda622411d8f868dff65c8fc95993463106fa09a3d1279a6510f760d18223bcd"
// synthesis attribute INIT_3A of bigblock1B is "256'hcd382b46840bab0d68f456dbd3d596c4d60080a853c78c7f58f548a21a230048"
// synthesis attribute INIT_3B of bigblock1B is "256'h17abb5e300006945014af24a51a8e7d613db0f953beac90c7d24a84e3db67e94"
// synthesis attribute INIT_3C of bigblock1B is "256'hcc0b966d71bb5167f6c496b8f9641edd2d98d6e435d5ba790710ba8868e81cec"
// synthesis attribute INIT_3D of bigblock1B is "256'hecce2ff4ad70f5b86956a029ae92106ddb173b9c24ec87798f382e553c2845f8"
// synthesis attribute INIT_3E of bigblock1B is "256'h2f4ff62e6210348ce817b4f316485de9c01020a36306509530dc32ab346be9e6"
// synthesis attribute INIT_3F of bigblock1B is "256'hc7ff012cdbd8cf2a81a6fd82a8cb5ebbd9f616a9362196d16db425424240e008"
// synthesis attribute INIT_00 of bigblock1C is "256'h2c6f8e5db656ad00190543657094f151c18302ab012f8e981f52c8589a39d5dc"
// synthesis attribute INIT_01 of bigblock1C is "256'hf12b089e53f11e98fc4d354e2624fa1885684dc70145580ce23c10bfff8ed20c"
// synthesis attribute INIT_02 of bigblock1C is "256'h4c61c51adf04441b582a8d2c5ee9054a000374f4fb720bffc322f2546b2bb2d7"
// synthesis attribute INIT_03 of bigblock1C is "256'he232ddfa8161562ad5b756e097d78dab49de9895149c6f749c907860a7a0137b"
// synthesis attribute INIT_04 of bigblock1C is "256'h809fd7f8cd5c411c9adfab577a060dd248f768b2c6da024880c145434c048248"
// synthesis attribute INIT_05 of bigblock1C is "256'h57576a8bc28ced115a6caf4e6c42e2a561410ec102c00e121dc093cf6183dabe"
// synthesis attribute INIT_06 of bigblock1C is "256'h672e446839ae754e151d817be2c9cd9a3deea77e9843fd354471a6b0a5384a33"
// synthesis attribute INIT_07 of bigblock1C is "256'h2d22b7123df236c2eda20ccc80218c5271b2d52f3561b1121c6607885e896a95"
// synthesis attribute INIT_08 of bigblock1C is "256'h764813d227022d6d1eac78a33fff00221400ccc03b0a5aa13f532f7b4047ef17"
// synthesis attribute INIT_09 of bigblock1C is "256'h9517eaba71d27aab926f402c2281ce57b853ff14f455b14f44609c67141c5ef8"
// synthesis attribute INIT_0A of bigblock1C is "256'hdf3b1267f6a102e77ef450097a50a177a71511ff5db6cf27808ebd8ef8b82b0b"
// synthesis attribute INIT_0B of bigblock1C is "256'h1e38a45ca6d2bd0bdf9ad71b793bd0cfdf523cfee6637f04f7bfd6433165f367"
// synthesis attribute INIT_0C of bigblock1C is "256'h584044a013750b952a28ad05439b18258f455d51533d800374f4fb7250ff1e51"
// synthesis attribute INIT_0D of bigblock1C is "256'h8308a9d46d13811b0021178cd6ca2976d777009ce347d235a113131caea88b0f"
// synthesis attribute INIT_0E of bigblock1C is "256'h0000993305d45569844bb1fae9c540201972f7d51682fbb7e6ad93274a8e0d2e"
// synthesis attribute INIT_0F of bigblock1C is "256'h78aba1fed6e94cf6ee8c0a7ddc604ab3ee5949f6a209548142f5d2f11a42a386"
// synthesis attribute INIT_10 of bigblock1C is "256'heed0247155a7522b53b38d022a9be043d86a47281ca35477528c7104bbff6d7d"
// synthesis attribute INIT_11 of bigblock1C is "256'h651a72e6750857f596b6408ad1bdb58152d6a81048eb0b3c8d357bd02a2bbb10"
// synthesis attribute INIT_12 of bigblock1C is "256'h56cd3277daa19c9aeff891bae3b94a0ec32e6a1fc6db2008c062a31f6592c5a5"
// synthesis attribute INIT_13 of bigblock1C is "256'he78d4ce3207efe65d49e84432c993007095831014cba561042afd8cf7ce6a01a"
// synthesis attribute INIT_14 of bigblock1C is "256'h9e32efb963145a558ecc5e931cd389cfdeeeb48a9ee0548c004803adc40135e7"
// synthesis attribute INIT_15 of bigblock1C is "256'hfb7219ff51d990f96599b9fcc6ed68f9b9ac4ad37f7ecea7c99e6c96078c3e82"
// synthesis attribute INIT_16 of bigblock1C is "256'h83156d9c900bd600c614df6c4c0425286c0da2bb302488165b312245000374f8"
// synthesis attribute INIT_17 of bigblock1C is "256'hd5661190e506db391b4a06591082a54031c62f6a1763ca67e147e74571e22830"
// synthesis attribute INIT_18 of bigblock1C is "256'h9e3a0092009c4588aea4460e2e99070d7f8c3b8a02bca3fc9647380932de25cb"
// synthesis attribute INIT_19 of bigblock1C is "256'he7fc74657436725378330c6bcf8c14013bc7f47bd45e0a236da37bc86a95e46a"
// synthesis attribute INIT_1A of bigblock1C is "256'h1c20ad4a50402c2f2441d27bc5251a04dd778ec6011892b2bb05599101a4583d"
// synthesis attribute INIT_1B of bigblock1C is "256'haf809e8c3d21e9f53e94fd0c6a5febfcede4163d09557d355a3851edf0b3e894"
// synthesis attribute INIT_1C of bigblock1C is "256'h0bd0dce3e0edd5fc717934b8b435aea5dc2425389634b49ddbbd463600414c04"
// synthesis attribute INIT_1D of bigblock1C is "256'hb399edcb323ffa8b9f0f9f72a7882aa8b70ac8c8a92484a624019122c4904856"
// synthesis attribute INIT_1E of bigblock1C is "256'hef9b6f2cb7da90cae0c8d8a6c138ccfca369d1a7e305a997ab4d477961cb56ce"
// synthesis attribute INIT_1F of bigblock1C is "256'h624b800374fcfb70e8fff30e2e704e9cdb72d7583d7557efbddf24ec9b0fa87b"
// synthesis attribute INIT_20 of bigblock1C is "256'h974d7904897e70a2ee689b0fd120231c09734c11e3889a2483db88262f45dcd1"
// synthesis attribute INIT_21 of bigblock1C is "256'h9fd7556e2bf6a89f63c836d81b6d2d030bc0f59014ad5a1270f5105e03cbe581"
// synthesis attribute INIT_22 of bigblock1C is "256'h2195044f002724b8514e0328e7a69d2838e749fc437675948417bf068bd79e1f"
// synthesis attribute INIT_23 of bigblock1C is "256'h6f460af305a643380fef38c37c3db2d2785a2839796d3f54ae09ae9a154c410a"
// synthesis attribute INIT_24 of bigblock1C is "256'heb529d0a69effab820907d293173ad15584a7af2868169a91f2d8e196523b7fe"
// synthesis attribute INIT_25 of bigblock1C is "256'ha36d59b50445ffafd6e504225656c7839d22877ce66dadd5e40e4c9faea3b232"
// synthesis attribute INIT_26 of bigblock1C is "256'h6e4c2405c4e4fd1c8d1331944f0a015f86d5a85444cba4ebb8d62f57a83cb2c4"
// synthesis attribute INIT_27 of bigblock1C is "256'h5594a86e07007cf70ae76b6abd0e6dd94d04690fd0211a68c00088511a092882"
// synthesis attribute INIT_28 of bigblock1C is "256'hcd7c409927a9d7ab2840a8f92c661b91646bc400f8786b7f197bff521b608c32"
// synthesis attribute INIT_29 of bigblock1C is "256'h25e3437849864b5c0339fa007274fffb4d3a4700b747391341df6377a79af7a6"
// synthesis attribute INIT_2A of bigblock1C is "256'h276ffa20fedff9fffeed5f0488b928250e2ec098ac7171a7a0f5580c25458b8d"
// synthesis attribute INIT_2B of bigblock1C is "256'h3daef6e0d62a58a70e80c4a6dd57198434988c1a20d1695ae8db4c296414d203"
// synthesis attribute INIT_2C of bigblock1C is "256'ha5612a982471eb196591249000b4114090249349ae55a4d6682a8a1d5fffb6a8"
// synthesis attribute INIT_2D of bigblock1C is "256'he34681e6a471989db0a47ffecfb7e94f99f3bdd7c9bb90f9f463058ac9b2e9ec"
// synthesis attribute INIT_2E of bigblock1C is "256'hb24a5af0f1649d33ed462103963f674a04cc243f3153c339d7adcba75652d006"
// synthesis attribute INIT_2F of bigblock1C is "256'h0c24657aa4ad6b6d0308e9b8711f41f46a42e3d9b045f0ca280acf06f7f26c6f"
// synthesis attribute INIT_30 of bigblock1C is "256'h8091ec1443502ea224ccebe853cc51c4f0a1756c19e9a83057a4a3a6886c9b19"
// synthesis attribute INIT_31 of bigblock1C is "256'h90243b9a7b1d3df407dd68f51ce99c13c44e699b8c657b2d2d4001f2801d1144"
// synthesis attribute INIT_32 of bigblock1C is "256'h54727deafbfe496420c832c95f11ed8546a7d4852d6e57d38b3ccff2fcf46286"
// synthesis attribute INIT_33 of bigblock1C is "256'h2e0b04e33baa26c417186988445d0330f9007274fffb92018b5c57d8e081f2e7"
// synthesis attribute INIT_34 of bigblock1C is "256'hd77f97fa33ba8715dcb98ef9a625911a4f6b1a18b45490ee60b09c5c75a48561"
// synthesis attribute INIT_35 of bigblock1C is "256'h3104ff54ad5f36f7ea11b597f916464e58a6fc5a4206c48b1fd68db58263a0e2"
// synthesis attribute INIT_36 of bigblock1C is "256'h2794ab12777fec5295d1233562cb3b89ede0b1c9e03458015151cc02ff29b58b"
// synthesis attribute INIT_37 of bigblock1C is "256'hbd553f42b4ac5e04733c0acb2284a3c24beb2aa336dc188ba97aaa3fc4f52666"
// synthesis attribute INIT_38 of bigblock1C is "256'h96cb3c5de9ba0ca80a31a465e5e331123082255dd9f5286f8fdd20c9da693071"
// synthesis attribute INIT_39 of bigblock1C is "256'h430d0643ee0e8c81db6b00d60001418088fe4a74f18f4fbdf76e3d975755e8ce"
// synthesis attribute INIT_3A of bigblock1C is "256'h22a28081d24cc1741733a199f048f0b80f775dd17ec3af35609979deda2bd484"
// synthesis attribute INIT_3B of bigblock1C is "256'h44ff789fb08d636362f0fd72aa3b876ca946b3419a6a5e6970942979055064e4"
// synthesis attribute INIT_3C of bigblock1C is "256'he83b259cbf55a1475ade8879aa981d43eabd6d15212f334837b178c8544f09d8"
// synthesis attribute INIT_3D of bigblock1C is "256'hac777124c929340b0d251b8a2a241f0851284adc033bf9807274fffb0bfdb7ae"
// synthesis attribute INIT_3E of bigblock1C is "256'hc0103e828fd9c6db024d40200030a3f4ffbbc13afa776cd499e01c6310ee2091"
// synthesis attribute INIT_3F of bigblock1C is "256'h0b68a821c79d628a1d0c18fe98a7563978c1c4d7017d2af4d85942d6340822b4"
// synthesis attribute INIT_00 of bigblock1D is "256'hfa42dffbd52c9fce2d63b0c272266cfacd7fab2e57bb60d0231400c2a301a0fc"
// synthesis attribute INIT_01 of bigblock1D is "256'heff3ad39242681629d7cf0b093c74181cf16116042a8115cd4252c9f58f446ab"
// synthesis attribute INIT_02 of bigblock1D is "256'h407294dda75b0b1e010aa66ffc8dbabfeed35e5177fb2ed5f62b4dda5c5c3021"
// synthesis attribute INIT_03 of bigblock1D is "256'h68ba9a90a004022f67fb3fd22f100629419292f499a26db6264d8a246108a306"
// synthesis attribute INIT_04 of bigblock1D is "256'h2eae8034b691424fa30e20f600148c4c14950f1019707a20a38afc28dab2a712"
// synthesis attribute INIT_05 of bigblock1D is "256'h86f6b6d79d22fc4054ef39b4b689dc085af1f50d26ae065c00e1fc14db40dd2a"
// synthesis attribute INIT_06 of bigblock1D is "256'hfffb83f9b3dc57ddfd167b5ed7f38e21af345cd9b9fe9555efe35550129b8bec"
// synthesis attribute INIT_07 of bigblock1D is "256'hf49390ed00b3a0576ee4752b880a20e63b7d2aa42e48c988595b0357fa807074"
// synthesis attribute INIT_08 of bigblock1D is "256'h6db4014b9515a6684bcfafbfffba9dafefffdc4b37e1dddc2ffbf117badd1518"
// synthesis attribute INIT_09 of bigblock1D is "256'h7dd7e94144f1185fc64847097d9476edf8e1141dbddb82ba26fd96332fd8be63"
// synthesis attribute INIT_0A of bigblock1D is "256'h624c95c76d49c400d5466d1364842ec1af3ab29c9023995bfa000b7315b4917d"
// synthesis attribute INIT_0B of bigblock1D is "256'hc7ad255ace64d00e35cfb0c3450322e697578633cc7c570c83a9eababe06e9b8"
// synthesis attribute INIT_0C of bigblock1D is "256'h1ccad128705eb1299d86d3f851295a9938ef430aaa378f5338a38c47c18c88aa"
// synthesis attribute INIT_0D of bigblock1D is "256'h5ea62e5f1f4feae8f1fc898625762a745b93ed522f04c3723968f3a267aa5555"
// synthesis attribute INIT_0E of bigblock1D is "256'haac4bdb346f6f58dbd3dfc7958d65b6bd62be3c3b3cf4ccd9b9555f0ec71d74d"
// synthesis attribute INIT_0F of bigblock1D is "256'hffacffffb81f4cfad6dfbf6e70ddbffff9ddc0cc69adffceff8ffd5bff5f977b"
// synthesis attribute INIT_10 of bigblock1D is "256'h1b44000374fafb7290ff4f1cff7c99a828d327d424920e531e61ce22b6a8ab9e"
// synthesis attribute INIT_11 of bigblock1D is "256'hca50615201a492702e6a9d0e8028548563734d09a37a9d2c241bc82bcc435cd0"
// synthesis attribute INIT_12 of bigblock1D is "256'h7b64d533484ac304072ac485c9545e8dd2d66ad1a00b21aaac2d01380bf22b1b"
// synthesis attribute INIT_13 of bigblock1D is "256'h38045b4370b0d0dedff16fa76ab8d7598b302260b88843242032b930dc2814f2"
// synthesis attribute INIT_14 of bigblock1D is "256'h608b20cd663b13289d35683371d83b12504995c040ce958a6720de622892989e"
// synthesis attribute INIT_15 of bigblock1D is "256'h6b1374a97ca6e29dbd58eb7a99c963fd96f66c531ba6f92df2d1597c3da1d225"
// synthesis attribute INIT_16 of bigblock1D is "256'hc9a8c1aeab011e3e263fe16672d8c6f025cdc02ed2310552e5d319d3ccdf2210"
// synthesis attribute INIT_17 of bigblock1D is "256'h5dab9d8563c8691bc2bcbc3a781bf18a301b1eeef17f6df5061abbea1d4eb169"
// synthesis attribute INIT_18 of bigblock1D is "256'hdd986c5acf03ad1e7fff597bb893e648f2b729ff0bf7d59a4961e59e89605875"
// synthesis attribute INIT_19 of bigblock1D is "256'h94cc9da42dda51a7d44f613098cc14fae1f77a9002ac50d57c25fd32ffffc0ff"
// synthesis attribute INIT_1A of bigblock1D is "256'h004661e05806cd64000574f6fb72aaff8db96665c210493452a8a5a96b2a06ab"
// synthesis attribute INIT_1B of bigblock1D is "256'h572cb13c35c648ad7b6400191ef02c0b030f8001199791601769bc0002c763cb"
// synthesis attribute INIT_1C of bigblock1D is "256'h46d01110cd6b19b9ddd504dadd826654f2522a7a90c00405796a7a802119299c"
// synthesis attribute INIT_1D of bigblock1D is "256'hb87d96e86d5223b8d4baa5668963e9ce4cfbd4191f6faddc0baf865c2478d75a"
// synthesis attribute INIT_1E of bigblock1D is "256'hf53a877ffed797847a84aff87efdd8342a1cffdf534cdd558e50eaab4c9ebf65"
// synthesis attribute INIT_1F of bigblock1D is "256'hdf0d820ef0f85f6f8e2048c286a9bae7aff40cea29145e00283f7de75bb18416"
// synthesis attribute INIT_20 of bigblock1D is "256'h55175f194a02b66261898babb62edd80e2d28b9d22229a8f8424f6d240544407"
// synthesis attribute INIT_21 of bigblock1D is "256'h96ffffcb04cecc8cb07f4c664e8ed2515042cdb76c4c4d5f738e58ca808cc456"
// synthesis attribute INIT_22 of bigblock1D is "256'hee0e265c25e824b7416b91b13aab6e6777befd4ab3663596b6cba346e2ba1e7a"
// synthesis attribute INIT_23 of bigblock1D is "256'h12296db2330a4945bac495411e5c84f5894c7b23afa9bffe95a673012c789d6a"
// synthesis attribute INIT_24 of bigblock1D is "256'ha000ace2422b0a192560dd4f1f3c00037483fb7257ff511119f677a332ebb92e"
// synthesis attribute INIT_25 of bigblock1D is "256'h5e533975f6f7315d8151a418f44f3497001b009c6ea45007710044ac33754c5d"
// synthesis attribute INIT_26 of bigblock1D is "256'h556a5e64bd97192e0d3d94cd2ba26a2ab80acb53d0f1f2957898a5327153a7c8"
// synthesis attribute INIT_27 of bigblock1D is "256'h3f299aed458fbac4d7bb64d8a90e5f6ed8ef9e5c51509021ccca988cef2a9eab"
// synthesis attribute INIT_28 of bigblock1D is "256'h5c468d37388ac79f05bd42382caa4a92e22e28a69b03f41e9f7fb49bd84d8aeb"
// synthesis attribute INIT_29 of bigblock1D is "256'h8dffbd2aa917b4413f4c6904415f2dedf7ccd608885a997a23724b6c8ace1049"
// synthesis attribute INIT_2A of bigblock1D is "256'ha302cc858ede278dc9b240f4ca74fb4f430f96c3243306e6e2c2d943bb9f21e1"
// synthesis attribute INIT_2B of bigblock1D is "256'hcd472d530194791fa5fbe915ae53fb313cb98e7f4fdc2beb6725b95a894b0ba6"
// synthesis attribute INIT_2C of bigblock1D is "256'h383a924a952411a3db940f413df7863bd0a959a8340edb4971b89224b069800e"
// synthesis attribute INIT_2D of bigblock1D is "256'h4dae120bed6b2caab3b540c7983159ddf6dede073e384bafacf65f57b6276dda"
// synthesis attribute INIT_2E of bigblock1D is "256'ha4a061794ced6724cc04423b4218851e5d692a4d00037494fb7066ffa766f573"
// synthesis attribute INIT_2F of bigblock1D is "256'h1a918085cf97f99ecfee43df3bc5f865bcbd83cb7db3d060310def3460887a68"
// synthesis attribute INIT_30 of bigblock1D is "256'hf70d24893e3658cc72541dffec0de9bb2566ef7d68f1c4eee96a548cce0d2993"
// synthesis attribute INIT_31 of bigblock1D is "256'h34813db82890a28b7f56958d240a4116ea47affe040748a3b5f38a77b8a7592f"
// synthesis attribute INIT_32 of bigblock1D is "256'hb56b3e4cc17016258f4bfec5b78973bc5f943d654c0890364dcb660d512a73a4"
// synthesis attribute INIT_33 of bigblock1D is "256'h629ad9362242fd2aaf79838133ab6ea598c6a2b4ff913b1dfa938bbf325f44fc"
// synthesis attribute INIT_34 of bigblock1D is "256'hd3bac7d4963dcb989018430a9198a9d26592a3b18a3ff4fab4cc9262232d8cbb"
// synthesis attribute INIT_35 of bigblock1D is "256'h0521aa412aa9c8891a0c545f13bdf6925f04880cb416e36d69a804885f7c460e"
// synthesis attribute INIT_36 of bigblock1D is "256'h1f71d012b3d0469fe73218cb23d28be64f72cb5457ebd34bdc49919180c21839"
// synthesis attribute INIT_37 of bigblock1D is "256'hfffbc6835dad88e871c31b2c3deeff2d13b4580e5792758e8d71c610291303c7"
// synthesis attribute INIT_38 of bigblock1D is "256'hf43106eec060947c77a4552b2c4c0cafdbbc18411792e9834add0351a0007274"
// synthesis attribute INIT_39 of bigblock1D is "256'h6b50596f356cd91c92e2df74871875752a75fe44b6bb209867392aabf2ce1990"
// synthesis attribute INIT_3A of bigblock1D is "256'h3a3ac12c34ad45de6ce031cec57ce504eea9411446db136e8414bb4817d82a1c"
// synthesis attribute INIT_3B of bigblock1D is "256'h8e459fdceb7404c90c45389d9bd1a5016b031736c71806b1099ec03724203a1a"
// synthesis attribute INIT_3C of bigblock1D is "256'h385cd4ee14eca1d98821afc85bb72cfd70141d7e587a60cae0585e6b620f1743"
// synthesis attribute INIT_3D of bigblock1D is "256'h924d3ff25bfff9fdce60d1e111f6f2d9f9fea85bfafbbebaad8eb992921252e6"
// synthesis attribute INIT_3E of bigblock1D is "256'h587a06e22200b845f491c521344a41f64a6b64a43691139212006d0298bf136d"
// synthesis attribute INIT_3F of bigblock1D is "256'h48b9b2f1903a27b1227bee9e13e4d7ce7addedbdc5ff55aa872ba35a8770dab5"
// synthesis attribute INIT_00 of bigblock1E is "256'hffe9fc735912a3048e8cb691313a61cc8c518d668d2a8584a9017a3e70b35974"
// synthesis attribute INIT_01 of bigblock1E is "256'h032cac807274fffb624b66d0e6cb1db2a1c12e90380832e18a674ea569a9342e"
// synthesis attribute INIT_02 of bigblock1E is "256'h08bfc11309406813846ee84b2d107343bd0d660c18a33b9d1ac21558e1884cdc"
// synthesis attribute INIT_03 of bigblock1E is "256'h9b67f9b6813c005d18044809908304652fe35682d1efba2f74c653cec4baffa3"
// synthesis attribute INIT_04 of bigblock1E is "256'h9e695d679bac58671090959f82546cc7c211162e6c976f7f6f1f381f5670b48d"
// synthesis attribute INIT_05 of bigblock1E is "256'h2fccfa7affb7c2cb65e74338f94e0cc820a7ac8e0bc72451538b754c85d2c763"
// synthesis attribute INIT_06 of bigblock1E is "256'hd7a072a87d5287d788803744300d9cc11b9f1cfb429250a1ee86fff9b387e660"
// synthesis attribute INIT_07 of bigblock1E is "256'h540716f58a7727cd2a170c0b29c80000001995a4a20d80deca97daa4cec3fb80"
// synthesis attribute INIT_08 of bigblock1E is "256'h60d336f8c6104911c039ed00689e02f5874351c328ceb890a14fde25a7280245"
// synthesis attribute INIT_09 of bigblock1E is "256'hdd3a7a1a67f4d5c77d75b39d59fe26215aa5d766e421459c3bda90431e95a395"
// synthesis attribute INIT_0A of bigblock1E is "256'h5137bc4e87db79290efa4a53b6d2098d92f04ed4d43e7a2bffb79676a924b1ca"
// synthesis attribute INIT_0B of bigblock1E is "256'h1e4849854a5c0302bb007274fffb8041009000006b803348d9dd001874892090"
// synthesis attribute INIT_0C of bigblock1E is "256'h114a9c18bb380e70d202b0782412876ea05a987471a78963260c04c33b8915e2"
// synthesis attribute INIT_0D of bigblock1E is "256'h6bfb2a9ca4cd23340c1a18ea50b76e9c42de56949ec6d93a9a2b1bb28724c835"
// synthesis attribute INIT_0E of bigblock1E is "256'h3bfef827653f418a65b48b43fdd52725d4e7aaf5c3b2d9a1729fb15a5382c468"
// synthesis attribute INIT_0F of bigblock1E is "256'h73a3a00851358b99b741ab98db690046a2c14735b1f4dca84bc379898612c257"
// synthesis attribute INIT_10 of bigblock1E is "256'hb596d1df6763956a662948da090b7c652140008180a8ea014d8df493ffacb303"
// synthesis attribute INIT_11 of bigblock1E is "256'h7eaf426424699efa3e0e9196ff01474e36ad552556a9bb503b33eab72d886179"
// synthesis attribute INIT_12 of bigblock1E is "256'h7a7da2f65aa8fd6ee46f5b74a857a2da67fbee953904b849498f7a499215aeee"
// synthesis attribute INIT_13 of bigblock1E is "256'h6012f0115cc02a12945f723b01907a1fd23a05c1d34941c60c24d7f81e579bf6"
// synthesis attribute INIT_14 of bigblock1E is "256'hfced6baf5134531cf1c5a8d5f172f10bc49f555c8ece6e95b925a291000aa800"
// synthesis attribute INIT_15 of bigblock1E is "256'h24291b471b62151051e659da0312cd807274fffb132cbccabc103190db667265"
// synthesis attribute INIT_16 of bigblock1E is "256'h26e0a7f7e47233f3792008029d9d845298911c34876dc066a44d69a718f5724c"
// synthesis attribute INIT_17 of bigblock1E is "256'hdddaf37f1fdf0df1f083fc781433c103167466c912c373c9393d22ff3353ca61"
// synthesis attribute INIT_18 of bigblock1E is "256'h01803c2a9ee90700b9df6b535b57cd4f8bdc6b38c14cffa605df907c3e00239e"
// synthesis attribute INIT_19 of bigblock1E is "256'h220e9e45162548c69a2b8d28592f1b5702c982cb3e09b844b100018101c55000"
// synthesis attribute INIT_1A of bigblock1E is "256'he2f50ef70b3840c2ee386c0f6c47b44a89c271294d4347a94bc9a0b23160821d"
// synthesis attribute INIT_1B of bigblock1E is "256'h0c71a2c70ddb1e956b0805d91ac2b1255d74c195c975a6905ea228ed69f37dc9"
// synthesis attribute INIT_1C of bigblock1E is "256'h0400b7547d73498346dc1ce614d9b64104e8404be50daace12ff3f84d22374d2"
// synthesis attribute INIT_1D of bigblock1E is "256'hec212efb28bfa7ff766eeb5f7246627134d5b895eb84a359a0ef9ba8463d0007"
// synthesis attribute INIT_1E of bigblock1E is "256'h747e57bba167add861149aecc8539d78910e3738bd487ed8add2287ea52b8d5d"
// synthesis attribute INIT_1F of bigblock1E is "256'h71a6810b264c04c7cb8a16e11638512858dc02e5dc807074fffbbf9fa576cbd3"
// synthesis attribute INIT_20 of bigblock1E is "256'h8fef0acefb39a9bd2da721957ed621f59422ff46911a2c99241607eee8662469"
// synthesis attribute INIT_21 of bigblock1E is "256'h0001801005011ca631bcb7f2e47342ac0333dad5058c98bca8e48fffa8565087"
// synthesis attribute INIT_22 of bigblock1E is "256'h415b8cd7eb7d2581028beb312a12e8a1720785dec2921ec0b85674fcc269c7d3"
// synthesis attribute INIT_23 of bigblock1E is "256'hdd1c0c67ac16a8b6dcd6472061ee9b5cb3b085263a50585c52d48c2ff2ab4969"
// synthesis attribute INIT_24 of bigblock1E is "256'h31c3ae96d59c472a8c36c7af09438a4d20eced08ea762b25c267bc3e810654ec"
// synthesis attribute INIT_25 of bigblock1E is "256'h32031197141a265131fadb4905460e80fff8ffffffffffffffff7fff20f46c8f"
// synthesis attribute INIT_26 of bigblock1E is "256'h5552e717b848791692b8117cfc4944a1000170060f2c8b3a170452ab86550954"
// synthesis attribute INIT_27 of bigblock1E is "256'h508847c3a70b0236d3e995c8834350ca172396addae216626e5cbeca3cbf950e"
// synthesis attribute INIT_28 of bigblock1E is "256'h2fff4623814652cc7362bb5b95849176fe3ad86655f55e4b22f7bdff6e48ff9b"
// synthesis attribute INIT_29 of bigblock1E is "256'had885b085ae8c60c776c4c4526806618021bb819232e5b493943800374eefb72"
// synthesis attribute INIT_2A of bigblock1E is "256'h07b0c5861039ab2e03fbb501f3be35502dafa9b1d228110977338551499f1498"
// synthesis attribute INIT_2B of bigblock1E is "256'h958a431e3ebca236181b0a1e000901004472b3b9b0b5df5f8166718ad3e8f28c"
// synthesis attribute INIT_2C of bigblock1E is "256'h591cf6e2fd42a48616b2ae1de36b352c242869b6cb837035c1dba15ac3be50fe"
// synthesis attribute INIT_2D of bigblock1E is "256'h35a19a8f94ead5ccb28d427da11ced84b0908ef52c48d3f478291040f838cd3a"
// synthesis attribute INIT_2E of bigblock1E is "256'h004e33c429cf56ca1ca10eabccc6dc396a85d81f2204e43ac67f65512d4b1aa6"
// synthesis attribute INIT_2F of bigblock1E is "256'h4716576d064e50000600d9cc2c49cf27c7dd95e24c61190f504964cf752848da"
// synthesis attribute INIT_30 of bigblock1E is "256'h3f71d38c8d919c5ffdb2b6c1c28de2d0ef1969c3d2d7ae0744714b4238c674ac"
// synthesis attribute INIT_31 of bigblock1E is "256'h9d6248b30219f0b55cc7662de704f485dbd21ee2d382eb5ac74f1c9bb34bfcae"
// synthesis attribute INIT_32 of bigblock1E is "256'h000374fdfb722eff75cdf26e8e50d15a5a6aa93c855d0b4475688be8ac9197d7"
// synthesis attribute INIT_33 of bigblock1E is "256'h2bbf317314986d586b8878a0c6180f6a4c95c2465a24e21b281c86165ac9a53d"
// synthesis attribute INIT_34 of bigblock1E is "256'h9c9e7b4cc6d37c9900f80b52a69c246d001781b0fd020bbdbf8e6501a9a64d98"
// synthesis attribute INIT_35 of bigblock1E is "256'h9fd1a1bbbf8a1d46b5ede84501de0126e3c40001014240e88743a1468da65f72"
// synthesis attribute INIT_36 of bigblock1E is "256'h72d97b96e1143d6451bc031e2435489e2b0f40d2b35d531fabeebee31b1f894b"
// synthesis attribute INIT_37 of bigblock1E is "256'h31ab2c432a1b65a9ed2edd31c4fc3c0fce69a447b5ae185ef88567efc7966f15"
// synthesis attribute INIT_38 of bigblock1E is "256'hffff3fff967ada96c79589f2ffe99adf0748abd589faf1a6a8ea6c84e583a979"
// synthesis attribute INIT_39 of bigblock1E is "256'h614913bb46d7d1655cc9b0be866c7ae70821b9076113b682dc918400ffffffff"
// synthesis attribute INIT_3A of bigblock1E is "256'h63e7d072c9e60d6e19ee5565a4b120239f973a19248e49260dceaaca80084bc2"
// synthesis attribute INIT_3B of bigblock1E is "256'hfc591034a9e8a91811e4ac41d16322bebce02fc89a52166515a18aebadae20cc"
// synthesis attribute INIT_3C of bigblock1E is "256'h89455b396a41800374fffb7242ff72a3a14e419996854db7d6548e230047a974"
// synthesis attribute INIT_3D of bigblock1E is "256'hbe1df6e16f8fff8239e314a06da87688fe20263c2f6d4e552810670c81db1818"
// synthesis attribute INIT_3E of bigblock1E is "256'h407c7e6155dccbbca33e64df58c1e115088344f968f038db00114080b33af21e"
// synthesis attribute INIT_3F of bigblock1E is "256'hbd37b4cbe29a92171dcb4207acc5169146fd138d6603e1b10501400031105c13"
// synthesis attribute INIT_00 of bigblock1F is "256'hf999d4326ef7dd711ef39c05b6f58eedd0ca67718ee644bd9e49ba979a3c8ff2"
// synthesis attribute INIT_01 of bigblock1F is "256'hb9105b31b4834184e747fd49b31479d4fd80dc8e22caca45cdd301d10d09dd87"
// synthesis attribute INIT_02 of bigblock1F is "256'hff02ffffffffffffffffffffffffffffffffffff74ff134f35ea1bd6ffc417ff"
// synthesis attribute INIT_03 of bigblock1F is "256'h005508003e705b282d80308e97303afee412cc243c3bf722e6a16da046e30000"
// synthesis attribute INIT_04 of bigblock1F is "256'h160c6e19bd248022fdbec615d31c951baac7f0197b92a578e79240b14e9b33f4"
// synthesis attribute INIT_05 of bigblock1F is "256'hee7c3fda026bee2133e42153e868356d963fc00e3a2fdb6af0b09b800f7521e9"
// synthesis attribute INIT_06 of bigblock1F is "256'h5708621b881d8b475ac1d14c800374fffb704fff3a99db04906da1236b382d46"
// synthesis attribute INIT_07 of bigblock1F is "256'hb3527dbb33f97fc6baa3877a58b6296414b06d687b077a80c6201b6a4bd9c912"
// synthesis attribute INIT_08 of bigblock1F is "256'h00235a0049c7cce905f33fcacafdd9e082a2338a694ab3dc5ad26d20b7244201"
// synthesis attribute INIT_09 of bigblock1F is "256'he09e71c382542ba340307a14d7450b06091ecb92e4451dd19812060c8a920000"
// synthesis attribute INIT_0A of bigblock1F is "256'ha079ea1ed5d557d9dbc86637344a7bc19a6c8aef72d298ffedd19a2aab1dcabb"
// synthesis attribute INIT_0B of bigblock1F is "256'h90b03488d5d8175eb69a67edd5fc70adb3cf5dd70fb53b165fd7c703775eb7c3"
// synthesis attribute INIT_0C of bigblock1F is "256'h957beac5e9d0b91b6d2a36e3e00cffffffffffff1d7facd5f7764faaa03c6dc8"
// synthesis attribute INIT_0D of bigblock1F is "256'h6e5121d9e3b4ca8e7b83596ddd0da22d0000a090c64c3acddca26616f98e8584"
// synthesis attribute INIT_0E of bigblock1F is "256'haa203b504d6388e9fa8b980c02939a56f0f37a0a5bb697ece4772df0c2b44ae6"
// synthesis attribute INIT_0F of bigblock1F is "256'h62460ffbe56e0e25fb7e85e3af8a9aa3a3669922b31a45ce8d8dbe96bd69eb59"
// synthesis attribute INIT_10 of bigblock1F is "256'h6cc61d310e4c05252b6a1c822f98318851db03e0ff807274fffbf6f534f45244"
// synthesis attribute INIT_11 of bigblock1F is "256'h2db99082f6b48d4e493c7750f4158ab792f05baf3db824289c13896d607220b5"
// synthesis attribute INIT_12 of bigblock1F is "256'h1a424a1249000602c60196010147a8d628276ea313c6794e030caa0b7d471b4d"
// synthesis attribute INIT_13 of bigblock1F is "256'hdf589430e506d0a12247d094af7d36ac8297269b01b9660e9901517c8d03c1a3"
// synthesis attribute INIT_14 of bigblock1F is "256'h6a3d4a22d91573f90bb59f9ac9e37d49c20893143d6154307e436ddb0857eff1"
// synthesis attribute INIT_15 of bigblock1F is "256'h56a02dad34a0f6df36f39c928824fe942dec3fd4bfdeffc2888bd4affd4891d1"
// synthesis attribute INIT_16 of bigblock1F is "256'ha820c580ff101f5db233de01975843ce15ca449a3342cb0b8997d35bb510f4ef"
// synthesis attribute INIT_17 of bigblock1F is "256'hba3182ee3ed8299b63da6ef15cc05bc82d2a2123f0e804d1bd851d5e5517241b"
// synthesis attribute INIT_18 of bigblock1F is "256'h91c4989813bb87c514077469bb6a239e324abbdf5c7ec8220835a42210b20d0b"
// synthesis attribute INIT_19 of bigblock1F is "256'h59f488d22eba29956e8963ef99bafeb92cbf74a215cd7457e1afcfaffe64df2c"
// synthesis attribute INIT_1A of bigblock1F is "256'h886d6069a0be6ac7892f064d05262b571a025d28c92f415a03abff807274fffb"
// synthesis attribute INIT_1B of bigblock1F is "256'heff576d06ef138b2380d3d9c947eb23600d88388f748099996f5e0bf1a015c81"
// synthesis attribute INIT_1C of bigblock1F is "256'h121c552e43473c15b08cc8c45e07db3e9ff88b7e1c50620ad58e880856079a6d"
// synthesis attribute INIT_1D of bigblock1F is "256'h676028b362825f2ae27f313470e3505c2f007252bc5149d4ddd925764014d645"
// synthesis attribute INIT_1E of bigblock1F is "256'hebcf5335e4dec76ed03be9a2b6c30b81ae72e91c49a9108a953ab50ee2ad6884"
// synthesis attribute INIT_1F of bigblock1F is "256'hdc7fc9ef3cec9a9aa746ade12d555c661a83c69180e123547b0ed3b79a95e31f"
// synthesis attribute INIT_20 of bigblock1F is "256'hbfdb9fd75b3545fe272a87280b23b4dc5fd850cb9e8c131c6b6ed3cb472df28a"
// synthesis attribute INIT_21 of bigblock1F is "256'h7b191daf67732de5672adab9b479729bef0d6398625d51b8bb7a30a5d61733b0"
// synthesis attribute INIT_22 of bigblock1F is "256'h8d7ece6552fd377bfffec6e76afd5ae5fabffa797dffd4cf79cfbfeeae65fd67"
// synthesis attribute INIT_23 of bigblock1F is "256'hff807274fffb579c189e8bd2944fc0c98d939e3ce212b585b6da1b6d92497e00"
// synthesis attribute INIT_24 of bigblock1F is "256'h2a068000ea9090ed00b7c5806fb4611d760d25063b772b042d58c9284bdb02d9"
// synthesis attribute INIT_25 of bigblock1F is "256'hdad9ade5230a1c6d4f58dceec5f23d891504136c9a508799501e1099325d75d3"
// synthesis attribute INIT_26 of bigblock1F is "256'h906b18ea817b5b42a5c2b6945a145f0d250a84a18a2d4cd5ee22a112393118e2"
// synthesis attribute INIT_27 of bigblock1F is "256'hd654518f06e55c171d707876618514435c781ec28b90805739466508eab0cace"
// synthesis attribute INIT_28 of bigblock1F is "256'h2daba05bf132827e88ce9ec2842e72c486ce37980b39a30eab73e1ec9e712cb2"
// synthesis attribute INIT_29 of bigblock1F is "256'hd7ae87ad798562df36c9097c1cfcaf376cc65f79e2e53e95245c14fb3386bcae"
// synthesis attribute INIT_2A of bigblock1F is "256'hb8846cde4689a41a571915e35b6a671e6833b9878d2c9cc3bd2fb9fb3da4696b"
// synthesis attribute INIT_2B of bigblock1F is "256'h1b6d924986008d65e6cb94a5ffe205f7eecbd24925a1fffe20cf2871d614c7bb"
// synthesis attribute INIT_2C of bigblock1F is "256'h06fe36661de1a83f29744b92702759d81747d230c18aa168d687ad7a01fcb6db"
// synthesis attribute INIT_2D of bigblock1F is "256'h066364580637fb007074fffbabe4e5788abc46b7692a257595d4dca245914a81"
// synthesis attribute INIT_2E of bigblock1F is "256'haba6940d584b31baf0000f1e8f2c010c8780601901910016c7bccb0346030000"
// synthesis attribute INIT_2F of bigblock1F is "256'h49b09e700d49d2a658d96e13abaf8f89dd5a9d71b68b29c604cad4340422d756"
// synthesis attribute INIT_30 of bigblock1F is "256'haf5afb7316ca51c9cbe58ff45ff2d7fb2ad67971b043a6eb3155acb49fbcba25"
// synthesis attribute INIT_31 of bigblock1F is "256'h3fdd5357ab4641a314f1dbe97c9fbf43bdeb54e8ff636c276d4ad0e3ff837f3f"
// synthesis attribute INIT_32 of bigblock1F is "256'h3295548c4e189052250bd5be1b070c257202936626db8f69c0912437f92134bf"
// synthesis attribute INIT_33 of bigblock1F is "256'h68a652a9d62bd499f3e69c45db5b5cb2b3f6d1f2eb849eacfae4b94e14aa797b"
// synthesis attribute INIT_34 of bigblock1F is "256'h91cac3476bec22ef094037a657fdae3c4f96402e3b3561976b5ef678b2bba32b"
// synthesis attribute INIT_35 of bigblock1F is "256'h325acb27b831f9e682f3cb7f45edfdf0482ffaa24d1699c8cc0d7a1111bdaefc"
// synthesis attribute INIT_36 of bigblock1F is "256'ha93ea22f40a1f46f2de1d12a7a390ee778392120e6f4b696e47148c0029311ec"
// synthesis attribute INIT_37 of bigblock1F is "256'hbae1e0eb0a1131205def222c80037485fb7220ff3147d1969249353604613413"
// synthesis attribute INIT_38 of bigblock1F is "256'h41dddbe7e4f6190ebd5351d2db4438ea0194eef4810d5aa8a6201b774d350000"
// synthesis attribute INIT_39 of bigblock1F is "256'hab0d9a61ceba77102437139440aa74d4e90f44b19d6d3d0784d3cdfd087bfd32"
// synthesis attribute INIT_3A of bigblock1F is "256'hac29efff9ff13939fe9d3e9cf87e9f08ba6d369495a7d167d8ec3e97d2734cfe"
// synthesis attribute INIT_3B of bigblock1F is "256'h6083f7fcafa84eb1acd03b29094436066af7391b185238026a1859b8c51bebd9"
// synthesis attribute INIT_3C of bigblock1F is "256'ha2a06552ab52461092807182dcf410dcea776282d24ead34928822683fa08a75"
// synthesis attribute INIT_3D of bigblock1F is "256'h5a252b5dfe9854f5705a1f80ee6aa05af2480a4f57b71245d5f354bc850961aa"
// synthesis attribute INIT_3E of bigblock1F is "256'hee7d233c1e56ea0b2a8fdac46cf5fabb3e16d2b72a0cb2bdd0f7ff1a17dff230"
// synthesis attribute INIT_3F of bigblock1F is "256'hcb46e8c13ba888d668a06f0835d19b1226b5d4c6b6931b8d1417a127c47590ba"
// synthesis translate_off
defparam bigblock0.INIT_00 = 256'h82ed003df1806b1c08610005c61c2b5f30a30400ee3e4eda04d604807274fffb;
defparam bigblock0.INIT_01 = 256'h7343a791b2859e3ca4a0811d1c98358b8a48bb10a602e15255c6061b00006b86;
defparam bigblock0.INIT_02 = 256'hf566d4be836d202b7f0868e1aaa89aa80cbebe541a80d1c3b949b60c8bc22354;
defparam bigblock0.INIT_03 = 256'hb84e1b5cf51ae993f3b60d185f24e93eb87ca8d0541234b3ab51a44a543ce398;
defparam bigblock0.INIT_04 = 256'ha2aace9a2a1be26f1d32e40d9a052b3abb9b89e5892426260ac664ccd523267c;
defparam bigblock0.INIT_05 = 256'h9ffe01dc140201c0c01ce57c34f151dc84267d447186f406ca444d66bacc28a0;
defparam bigblock0.INIT_06 = 256'he79e148a21bf04401d257933edc12b4fea720674d632db4783036db2b6dbdb6d;
defparam bigblock0.INIT_07 = 256'hc5d713590184c7bfef7c1aa3cc78df40baf1e3050af10400e0001b07c68896f3;
defparam bigblock0.INIT_08 = 256'h905bbd0b114c84e65f786d83492400ee40000fe91b4160c62385b3e1cc88e8e1;
defparam bigblock0.INIT_09 = 256'h0e007274fffb3722907f6cc6445ca899bf8722cc40e4a32b012770ab4a2e9020;
defparam bigblock0.INIT_0A = 256'h7ad18c11245184ae2848a0db71a4755b304f0c42cb8a126040785126265c02d7;
defparam bigblock0.INIT_0B = 256'h705dbbd521040940a090e631d5ece5d45154753152a13bc5b5cf420882972699;
defparam bigblock0.INIT_0C = 256'hb05cfe22fd48c4197d88392639acb1747904b410a308d1e06cd8b84e516d8932;
defparam bigblock0.INIT_0D = 256'h8a9b680872238b809b8300000a20002336c2fc71d4ad8410c3abc4f424889249;
defparam bigblock0.INIT_0E = 256'h6cefbe2d95dca5e43892acbdf1ac4cc19131c3679e24411bb520d054031884b9;
defparam bigblock0.INIT_0F = 256'h162e8b0ad12faeb96aaa9289b48e44679b6a974ad2afb65844bcd8fa4abd58cb;
defparam bigblock0.INIT_10 = 256'h487b0802cbc12922e3cf1689284362d3047263389b907e824398345c58a55848;
defparam bigblock0.INIT_11 = 256'hd9233341fe6a0b51159164cc4350852cffff463fc840dad9e19c2468914bc2a6;
defparam bigblock0.INIT_12 = 256'h6b68fae5b36e28e476c2037ba45922832115a20a03074078330c4e47502951a6;
defparam bigblock0.INIT_13 = 256'he92359de03381b807274fffb6fe9ddcdaa5d94b39988da759665dc291939462c;
defparam bigblock0.INIT_14 = 256'h4c86337b846bc9088c81741407efe07198697ba44947120c0502bbdc17812dc8;
defparam bigblock0.INIT_15 = 256'h6665cace8eedea3163191e46fee4a18ecf621a543151373ba1462d74c2d11851;
defparam bigblock0.INIT_16 = 256'h08d48a39c1018f26409aeecd17403304fb05bfffdb4921d2663b69abc99cb95d;
defparam bigblock0.INIT_17 = 256'he418922d95e48918bb6f48fe6d02d178708107e437a110b70ba8448294d40c44;
defparam bigblock0.INIT_18 = 256'h41c24629de98ce6705faca792891bbcab320456b3952d126a1fa0516114d04ad;
defparam bigblock0.INIT_19 = 256'hf0850b2a71545841462ae67af485690bee5e6dd75e12b5943274f87f3cf75c05;
defparam bigblock0.INIT_1A = 256'h2410890ca1438f0f07809a338f2f7822344859dccf30b6d9e36d6536010049a4;
defparam bigblock0.INIT_1B = 256'h5c223b4d4fbc3ccb892c962d9761c0eb98d2e2945683a8acdba83b683a004b6a;
defparam bigblock0.INIT_1C = 256'h3ea37bff379dad7d489154af964f1b91c63a36fcfdf8cd2531f2d39b168ff1c8;
defparam bigblock0.INIT_1D = 256'h9bca18021e48612648de032528007074fffbed47f1a76c296f961dfed422357a;
defparam bigblock0.INIT_1E = 256'hf174e233cabd6431dff6b7d60c9d8468241104efe059187178c3651b344b0462;
defparam bigblock0.INIT_1F = 256'hc21187e6ee9515f9ab9182a55ca198ab781a6d86b91bb2a9fc00b52b5d513114;
defparam bigblock0.INIT_20 = 256'he7efb2ab5acaf870ca6563460de818df8b4b74aed864736ec414f9d23c48a100;
defparam bigblock0.INIT_21 = 256'h854c14686ea1956e3be58a2db0a65e1b12e5927128b9bd101a9dbb33f9add8c1;
defparam bigblock0.INIT_22 = 256'hff261bff400890a405089fe41e55c18b8806174e2c11cbcbb87d653253d7e320;
defparam bigblock0.INIT_23 = 256'h056f84df32213f440916008b2d809901ca994f892c8b86872575732ade9b9f01;
defparam bigblock0.INIT_24 = 256'hb79d63def3842c7d87cc71f2f8cf66ceef633b6895658e3964d0dc9033cf234d;
defparam bigblock0.INIT_25 = 256'hc4a45ce785c569b2768f9b82c2874143ac44309496b276e09db92738d079f197;
defparam bigblock0.INIT_26 = 256'h40130100d680d3a9c19c23db60d2b162a38112937fe6afa9f78d2fb28d92cec4;
defparam bigblock0.INIT_27 = 256'hfd774b040302bc04a13b881623375dc95c488003743bfb72f3ffe92c92567fff;
defparam bigblock0.INIT_28 = 256'h2489e82f000254c9e801be00d33a6d5eb7d524bf0808200c2ee44f0567c04498;
defparam bigblock0.INIT_29 = 256'h74e7c10e8935c1f18149eb2c5b24b2b4b8d94e35d21001f08c83e0b667971a4a;
defparam bigblock0.INIT_2A = 256'h1e26a6bc508d15ceff21e949d8f3ff3ca23bdd56a4dfec21752cd0489a9e9d48;
defparam bigblock0.INIT_2B = 256'h133db1edc6edeb9ca446ee8cfff041afe0116b622f3e73cdca637f8303d02506;
defparam bigblock0.INIT_2C = 256'h6a1b3aefa9eec57948baad41412213a285642a1012a700293640094926ba6a94;
defparam bigblock0.INIT_2D = 256'hd7bb90020f95fff7289e7ceb437dcbec3ccc518e8655912ac6c44e2b674ee8a9;
defparam bigblock0.INIT_2E = 256'h9bba472274ab0b34ca0313d01505b4bb2dab8cf5219ebba0885d14a8d699cc14;
defparam bigblock0.INIT_2F = 256'h04d3c151b8c67dfbb677b5a1cb7144ac3896b1a0d69abffe10414a406ea85073;
defparam bigblock0.INIT_30 = 256'h0c529c45297bd08ad265c8fc2709a5f8b0adacf510d7844d89a3b4d3012a0990;
defparam bigblock0.INIT_31 = 256'h67046f40a62427754c612340ac20a13bb0188615dd690d3f8003744ffb7204ff;
defparam bigblock0.INIT_32 = 256'hd6ab523fa91fe1458f0a9e604770ffbfe4c42efeab66841181bc803d348ceeb0;
defparam bigblock0.INIT_33 = 256'h0db1f5ec8e6511dbd965df4ce5eecd6154a4174fdab71d4da4fa6998ebd3655c;
defparam bigblock0.INIT_34 = 256'hb25d6801660854d18c1f54a4e58ba7610a01d41108cafffe892b5510a6401ba2;
defparam bigblock0.INIT_35 = 256'ha926045523efba904f18c3e6af0a222daa35bc8c2aaea2a1a9652ead00fc0cc8;
defparam bigblock0.INIT_36 = 256'h5feee7fa5e4e2a8e11c862a338bc0b29f4af27df9efb43fdfc67c4ebfc98295b;
defparam bigblock0.INIT_37 = 256'h2be097f6d4718696c01909301532973820f6718bc82ce2a15652a1b181f2db30;
defparam bigblock0.INIT_38 = 256'h1520080088b33a017ca470e846d128bb7e5d7e87c3391c290e48b0c26fffa046;
defparam bigblock0.INIT_39 = 256'h85d25ea30f6d8b7f1637f797303b12936c2cb890e28962e997700e2a9dcd4399;
defparam bigblock0.INIT_3A = 256'h745ffb724cff06ce3b424d2e00e4cf0661558412a8e121d1534ff3bac0b4242c;
defparam bigblock0.INIT_3B = 256'h810c248c6ea46d0a6bc0a7a403754c6d2374a90c229ba01887335d6112340003;
defparam bigblock0.INIT_3C = 256'h491e90ce925a8600b7ae6e48aa8a4674c0ddececfb76a7fe934ef334e558da48;
defparam bigblock0.INIT_3D = 256'hd24042526554a3ea02c251aabe9585317cf5dc0caa6215cc9c660f56fffb1d4a;
defparam bigblock0.INIT_3E = 256'hd38da0a85736af35ad8990c851f0d1bdacb6ea637b15b42e8dc833551f2c014b;
defparam bigblock0.INIT_3F = 256'hab322b6ff3dd673bd7d092a22c7d2b5190bada40d56bd5552235846682acec2e;
defparam bigblock1.INIT_00 = 256'hd634e6c7fffd24b7851860596b569dec774a40f88300ef4347b1c2c156540d7b;
defparam bigblock1.INIT_01 = 256'h2c91b674a9c82995001ab1f010128a4038ad20b1213b0625931f163c5369b1d3;
defparam bigblock1.INIT_02 = 256'hcc7a42bec111bce5819863ca6c2887a865cdd8ca134f6c63c88ce4415cb0be1b;
defparam bigblock1.INIT_03 = 256'h8b46377e05c3667171d0d191c1aa09b03eae9909d631c458b324813040626184;
defparam bigblock1.INIT_04 = 256'h5e69de3d8002746dfb7000ffa0396be176f168d57533cc38a30e2b9f3599a544;
defparam bigblock1.INIT_05 = 256'h6db226db1272980013156f34758a6d2083241f794c552234cc18429bf01be929;
defparam bigblock1.INIT_06 = 256'hb02918578000713a8464cb284619c07349483dfade067e0b94bf078647a919e4;
defparam bigblock1.INIT_07 = 256'hfbfbf71b90ead3596f45c73e46d15354df0facf50871307aac363094d56aa2ec;
defparam bigblock1.INIT_08 = 256'hb2acb7470523eee2dce88569e32ea33534a24e3dc5a528e1a63851ece7cc14de;
defparam bigblock1.INIT_09 = 256'hd9886db6c76b022cfda09ad7a6b510265f2c60aa3053a170203af9272d63b7ba;
defparam bigblock1.INIT_0A = 256'h50a641bb51390001e471282c96924e33427b8d2b85165cdb3958e0c27a5287ba;
defparam bigblock1.INIT_0B = 256'hec5bc25bd76b24a323d81ef0be4ca4d191fde706acab903f0483488675639dd7;
defparam bigblock1.INIT_0C = 256'h3e8aa8c62dad0efce5b6b265778fba515cd4dc11983339f160b70ab447d79cf6;
defparam bigblock1.INIT_0D = 256'h25e5a2b5c3cddb6c55b638ed40682cd01eb3886138d85010f87c0ea488964583;
defparam bigblock1.INIT_0E = 256'hdbed1c222b6868c9445f030e7c807274fffb409e1cc50472284c4388c13d0b21;
defparam bigblock1.INIT_0F = 256'hf654cf8138b2880551b4121345320d49b41389ef6074a46f7da5e10f740b0826;
defparam bigblock1.INIT_10 = 256'hc0d19dfd6306c730f3a3fb5392c9ab4cd8a4d627c36031605ae58af098a21718;
defparam bigblock1.INIT_11 = 256'h68d76d697b5dd6e8b96eb6034a9e1fe8c76ac49656d116e5b50f6ed477ddcbcb;
defparam bigblock1.INIT_12 = 256'ha106dc22a6e62e8efab257ff094e2a04b4ff5aeb7eae0397820d5705a8517335;
defparam bigblock1.INIT_13 = 256'h91691f79d2cdeeb931f13469222d033eaf00ae3dbf13c5c1b2160110c813be82;
defparam bigblock1.INIT_14 = 256'h9214fdedf682fe8bfc881f75834558c20e19a745ce21fa15f5a77ec0284ca4b3;
defparam bigblock1.INIT_15 = 256'h255936fc7e6bcab1b37e8f7da23f6f0ff3f09e5e25216a9d75ba0c5944f8c76d;
defparam bigblock1.INIT_16 = 256'h8f8006b54de169a4b441fe5197ff82828124a14421dd2d94815a65b8ebf8bde1;
defparam bigblock1.INIT_17 = 256'he0c824fc1f9c04cd61f397001c89a865000004048ad0846535e9f19f2bc69049;
defparam bigblock1.INIT_18 = 256'h511d704c0c43fbbc1bc11450e986485d02e88a807274fffb2fe77864e0e6b69a;
defparam bigblock1.INIT_19 = 256'h5fb8ebb189ccfa673dfcca67a27d1c031f24f58e0d88f0110b6ea06b20d67726;
defparam bigblock1.INIT_1A = 256'hde500786148436cb9355da9da7b1820e6e5c9af9fb9d3ba95d667ceb3606363a;
defparam bigblock1.INIT_1B = 256'he55e9065d96315400437d4a3b1625fff390133f7e755bbde1322d1020b35030b;
defparam bigblock1.INIT_1C = 256'hf363e0ca60cbc68e32afc1a625857a240297600083115a40c30077c6909a285e;
defparam bigblock1.INIT_1D = 256'h7c4eed36923b957637fb6e5c6cf7563103e5a66524864d3a2fb9e292f152928a;
defparam bigblock1.INIT_1E = 256'hca315e6d4404596cf044b90f335c9c5b7ac6bb71c36f8840ee3910e67dfc1582;
defparam bigblock1.INIT_1F = 256'h8eca8dcc0996e0ab305868613695fff8221700b3b6313c584b182753f9cc787e;
defparam bigblock1.INIT_20 = 256'h20cce2f524e02023fc78842c9a8d0220469ad1518000997684897647b50933fa;
defparam bigblock1.INIT_21 = 256'h61de52d865b498abb432ef719b52d6d7bc5572a285d1529e7836221b2029eac3;
defparam bigblock1.INIT_22 = 256'hc06a246d71a69cf9604c0c25db891a4114606926415c03029a807274fffb61f0;
defparam bigblock1.INIT_23 = 256'h42d8beb8b3ba99e8d5a18faa9da4d07dcb928da3fa5a5cc9f35c883024218b6e;
defparam bigblock1.INIT_24 = 256'h5a745839e496c640f68f95ff22e427fc21d4cd8b4282b69d52e709be4a1d3450;
defparam bigblock1.INIT_25 = 256'h8822848253729d3e4ebbbca9026f741e0013a24d00222d0975cb1a2a4596f49f;
defparam bigblock1.INIT_26 = 256'h718ff7e9d0a0651fa53dd8a6a7ff27127cc22291c438c1a4ebb1900fda8fe263;
defparam bigblock1.INIT_27 = 256'hb9439be6f02972a37f4e41272aa253042659f48d84a549923f2d4fcfc96731fc;
defparam bigblock1.INIT_28 = 256'hb3a82e458f767e81e7da428289da52b3f65545ff8828e8ac575fe292faefdcad;
defparam bigblock1.INIT_29 = 256'h542289ab71093fc119e43a7be624109384678b395c23d3c6cf33000019104728;
defparam bigblock1.INIT_2A = 256'h69dc9d5504139ea93cba6b884969b8cb4953aa199efcc9301024536afb1716e5;
defparam bigblock1.INIT_2B = 256'h7074fffbee4551b585416135a5ed82e42ed4e2abc903ceb86c05c0ec45db6d7d;
defparam bigblock1.INIT_2C = 256'h88c9a460872ec859987275a41925500c0c43dba91741430848c7445d0335a880;
defparam bigblock1.INIT_2D = 256'ha6ad70c4eb73632907c88957000fee8bbb92e34d00060600f68fc6ac12602fa8;
defparam bigblock1.INIT_2E = 256'h7367d23c5bf77328355c3301d86ba88d2953240dcfdc655d000b000554395244;
defparam bigblock1.INIT_2F = 256'h8bf0d7c2e396885b7673bbba2c29cbfe1f0a5be0699d126a8fb0a24b72156069;
defparam bigblock1.INIT_30 = 256'h5438ba7b2ab44abafc075e4f3ffab9d4eafa3f3343bf270f8b29e29d07c6b6d2;
defparam bigblock1.INIT_31 = 256'h480500c0cbea2b8ed7309f45a2338272fe9a72a8682e17cefbf5015f10a0ad3a;
defparam bigblock1.INIT_32 = 256'hda00d8194a566b9e16b2938c3cf5377e48683aeeca9ae17650f767b33f1a7880;
defparam bigblock1.INIT_33 = 256'h1f5346dfa50b90a35842dfd60bae49063e3e482b453673d6cdf0cc862a2907ef;
defparam bigblock1.INIT_34 = 256'h04044040ff019574d259dc592abe9b5436bc25676154225435480f552892b2c7;
defparam bigblock1.INIT_35 = 256'h5bd12034800374b8fb72c7ff67f4f74008caee9a68dd2151302caad22611e36d;
defparam bigblock1.INIT_36 = 256'h9002c18543c94934360c6de4670775002618276f0bf1653a7a18c29bf01a8941;
defparam bigblock1.INIT_37 = 256'h93908b662e0ff49d62d480cf7291b4332a1c1ec6212c5035e52258f5000a4480;
defparam bigblock1.INIT_38 = 256'hef3d052e4c8c36e12a5bf0a5eb432cd3bde4635dfe0c372ff689d0dfffc42b6d;
defparam bigblock1.INIT_39 = 256'h031ca59edf36694b9deec570042afced2edaaaab3222423122d26e6b998e7881;
defparam bigblock1.INIT_3A = 256'h4ad85626a2252f9208c2cdae4945815ac55c81f3d0902547fffc002b8114c5c0;
defparam bigblock1.INIT_3B = 256'hf2290fe0e1cb74ec6467c5bcc5a84064aed4b3d524986ea975a0dccf2025d549;
defparam bigblock1.INIT_3C = 256'hab1c227790a3c0a726d5c8e0d07c8ab64a8cb91ae8320ae58197b1f363e6bd30;
defparam bigblock1.INIT_3D = 256'hed47081da1ced33e8e36985ae675908639b6ed12a9ee805df749a41674dba690;
defparam bigblock1.INIT_3E = 256'h1c92319998516b69120de886615e347f74f18465b54e91d5a33fa8aa20f6cd55;
defparam bigblock1.INIT_3F = 256'h429bb01d862d5be1f838800274c7fb722cffb389e997db0826ad4dc98a8d9202;
defparam bigblock2.INIT_00 = 256'h404d518fdf73e8456b301bee20d414886df073095880a620316f4ca125167d0d;
defparam bigblock2.INIT_01 = 256'hf925480a11f071212544ed160948066a1411043bb0944a3258c8226391ff3e54;
defparam bigblock2.INIT_02 = 256'h367d200c5a68fda41e31d4f0c4cd5505125047f11aa2c8072385883a63069f17;
defparam bigblock2.INIT_03 = 256'hcddfe9bc14a7be3bd9f5539c4053dd158b6ce9ba43f68f7839be5429b5951b69;
defparam bigblock2.INIT_04 = 256'h7eed77b6ce4b4c85d434d12953ab4572248b68b08818cd81b329b5cba6d0956d;
defparam bigblock2.INIT_05 = 256'hd36c1b7be3a86b2f55203c469e3433badee6ce8d528b157e64e7e9ec99a5cb1f;
defparam bigblock2.INIT_06 = 256'h8d7db514c82d0ebc0f91ad2aea0b2df44a96098d6717659182815525eaa0bca9;
defparam bigblock2.INIT_07 = 256'h55ae946d5bfdf6a12cb9bd851864babc3aff23211876563e377620b124cd2b4d;
defparam bigblock2.INIT_08 = 256'h9fe9f2d22f79cf9e6152de2c55d38bd55b5a21120979d10219ad098e3bb47169;
defparam bigblock2.INIT_09 = 256'h4b78c208dd0464bb20296615ddd19929800274d3fb72a9ff967b560e4b2faef3;
defparam bigblock2.INIT_0A = 256'hba3e86f46c235991b51f5fa75859fd277f5a394651192ff49b106be0a4a4937b;
defparam bigblock2.INIT_0B = 256'h9d13b2c74a1793c21292c2850680e2af87a9c3a55dfa30089ae1482a0219d51e;
defparam bigblock2.INIT_0C = 256'hf2526cb2b074455ce3eaad363dee1c9a9ee5b03bb492e56d50a6009327b41b75;
defparam bigblock2.INIT_0D = 256'hd0459a6dafb8f2599dbdc5cb98589ce07b2a9e655e386c09002e420019550340;
defparam bigblock2.INIT_0E = 256'h35652af14068648fee4a4b90eeea0c33cddc4b132c213121495075143ba6ba99;
defparam bigblock2.INIT_0F = 256'h5b9590ba32fbe1022a95b492a297e1c077089d1ae06b36965af804c4cebf43dc;
defparam bigblock2.INIT_10 = 256'h994ca740440a1ec89389d5e3fffd23decde16904f5321ec6907f17981e0f1056;
defparam bigblock2.INIT_11 = 256'hc8d2a5c2d1d72c4b9fe7c15aa52a0b20a6250410eb28c285782350fcd47fd118;
defparam bigblock2.INIT_12 = 256'h2fad69afc9a6d096dc79faf718c54ee6fa2fcb79e1e1dee5a3a0233c51cc4a28;
defparam bigblock2.INIT_13 = 256'h7120a430a77f4b9402b2fd09e49b4028cc2c5ee8cd29000274dffb707bffada6;
defparam bigblock2.INIT_14 = 256'hebc54a78125d0185cd09e500c985138c3e08ecdd16adc6777ac9011870f4738b;
defparam bigblock2.INIT_15 = 256'h58b8564363a628084a7546d25852211a2e02b308b810a163ee8269e9c3af05c6;
defparam bigblock2.INIT_16 = 256'h9be6e1db355f2f2b9718000798405e2920a0da82b3d53c48bd2415cccfb31c63;
defparam bigblock2.INIT_17 = 256'ha5c2e750259fa4ad5b0889444798b6d4ba86302a18f32f93a069488a2ab4a7cb;
defparam bigblock2.INIT_18 = 256'h2cc9995d2f46ec55ff96274962b7591b5e375c93b5fe46ba2aa87b9c2cb6b6ef;
defparam bigblock2.INIT_19 = 256'h8dfe66cc22c1404d6151aa2e54dc25a31b6b67efe63eebec1c439328abeccaae;
defparam bigblock2.INIT_1A = 256'h50c62f149c77e174ec81b1cb903404f0da4aa1990c18e617db6811b60c1c8020;
defparam bigblock2.INIT_1B = 256'h71f8256359de3bc663baa97db3b6df7608740a127e34cb84912971d8420ad842;
defparam bigblock2.INIT_1C = 256'h7274fffb297cb6afb5cc985667a57a6e36f0d4e6cc48c858dc6c3f2af1327d0a;
defparam bigblock2.INIT_1D = 256'h8d88b4348b6e807c185175a6f0c9304b0c239ba91c021e4a512851dd0373eb80;
defparam bigblock2.INIT_1E = 256'h496deb3a0aa016275bf7ee55ee5421bfe46d929f74c5c4547a9588dd707f7dc5;
defparam bigblock2.INIT_1F = 256'hbaf314874d5086f4c28306286952391b3cb24058dfd8b30e6e3e3d4d1a7b3bbe;
defparam bigblock2.INIT_20 = 256'h6332c93f509462825cb6f71b29246cabc17507c55800000890eb0092a7b57ce6;
defparam bigblock2.INIT_21 = 256'h5c50121f14384af34b75c3901b7ec4191a9fcd223f4ebd04f8132e32fdac879a;
defparam bigblock2.INIT_22 = 256'h5b1d46fb569b6593ecfd9f4ad4f2a9c66cc822e6de84d86063e259875dfaa548;
defparam bigblock2.INIT_23 = 256'hcc6f44c72187946c71b410838280fd5fb3e250e8d72e25020ab75044050203c2;
defparam bigblock2.INIT_24 = 256'h91bb6610eba91e9a8349f681e00020520200c8888856f3a1541d883aa1b45ac0;
defparam bigblock2.INIT_25 = 256'hdc726da6caf75631c15af5b4c3a708da7e02bf2804be248264d2e0986ba39c16;
defparam bigblock2.INIT_26 = 256'h4d5c038ff2007274fffb951373bddcc833fd9a4d5b3558e45b2882107b7bae60;
defparam bigblock2.INIT_27 = 256'hfa2921a4f523a0d16830876e0871bd6d73a4f4cb604c0d889b9d21221cf8e9e9;
defparam bigblock2.INIT_28 = 256'hf690cf19ed39f09f77fd48699bdd7de0059c5ce763b55ce354ddf8c5d9be8910;
defparam bigblock2.INIT_29 = 256'h012b589a549265246410519b19e56a831ab38074b9a88266c3c1a490dc6d41a4;
defparam bigblock2.INIT_2A = 256'h9dd066071215065c201ebbc9e0ec16f1a54fa3bdc586028e8f3db64c4da14387;
defparam bigblock2.INIT_2B = 256'haf0c79cf6f931fde5a759ebe37fde3ee089dd8de479c8ca1a379f943c5cf6849;
defparam bigblock2.INIT_2C = 256'hb6db9cb80136f214b8ca6e48a13b8d2a3a3c042a3a093e3cd2482e69890cb58b;
defparam bigblock2.INIT_2D = 256'hf48cdf87f39f4e6848ba0808b3c9d169ff79f815ce7708d1b0a4908f2a0754a2;
defparam bigblock2.INIT_2E = 256'ha77471e9e6b7fd7aa13f3690236a86db64d822db00295b1a9a7f68a87bb1941e;
defparam bigblock2.INIT_2F = 256'hece597dceddc472ba84d4b3386586443688a8a1be5acd2fceec699834c12b9f8;
defparam bigblock2.INIT_30 = 256'h1ba24508b12c475b0349f1807274fffb13b9849fd24e90405385e2f1274c6a09;
defparam bigblock2.INIT_31 = 256'h80cce8d6b4581e848d8ef9a294d0dc200a6da861987c6f84c125740d18a33b7a;
defparam bigblock2.INIT_32 = 256'he872e380fd1df29240825a15f567b4951b8d465942d2b34ce87ec99122279320;
defparam bigblock2.INIT_33 = 256'h46acad8ad365054eb4485c7111048726cb7abcbeb7b60e5e273585ecf23ce8aa;
defparam bigblock2.INIT_34 = 256'hbe7acbdaf55898f6e007e95198c0e064b4b8fa18493765bb88f330b2639f5ce4;
defparam bigblock2.INIT_35 = 256'h895835262153b8ed352f7dee26f7cd4431db97131e943b8774f1ac7dbbaa251f;
defparam bigblock2.INIT_36 = 256'hcd67af2ab492d38d2108fc01a5499d8aee49f88502711830660d4f2aaa7eaba7;
defparam bigblock2.INIT_37 = 256'hcb9b68e51664c201ae7c949952dca247e65e46b84f33606b52cbfaaf1857457a;
defparam bigblock2.INIT_38 = 256'h2db59dca041a7b38f2ec5327e06c0640b567ed39609580588aa15544a94a7d56;
defparam bigblock2.INIT_39 = 256'h724ba11781357ccaa14bdb1e3ae191dea2b5ee9b599ccbef7c435d24b61393a9;
defparam bigblock2.INIT_3A = 256'h604c0cc3abbd2b841d28e96845dd0304f7007074fffb58f31200d131896e6196;
defparam bigblock2.INIT_3B = 256'heae853985ef644b380c0754119480c25e0479d08f43092eea0a6a45677a72ca9;
defparam bigblock2.INIT_3C = 256'hb1008bac0e9b3951e8c91e758dade40132f5297029e56233b7d9db6d5cc65504;
defparam bigblock2.INIT_3D = 256'heb8dcdcbde6109a4e16d6add178b110011b714da2b200b4af49878ea1aa6f9e6;
defparam bigblock2.INIT_3E = 256'hcd99e4f5a52fae6c512d1d06719cf554dbea0ec744aab3bfc567f7cfa4f791fd;
defparam bigblock2.INIT_3F = 256'h60cb2eea68f732ecd4df14382dcaa16ea73d48a8618bcc88b5df79e27149022f;
defparam bigblock3.INIT_00 = 256'h91e5346d6d83b51b49298a264720cfe8859ee173d9c0aaf8e879d1ed86fa14f4;
defparam bigblock3.INIT_01 = 256'h0679b003675024ecda2b127e7b4a18cfb0c0a752a15e75a9e022abd4021fbd6d;
defparam bigblock3.INIT_02 = 256'h4b3b9652452c9e9127222f6e76c5285464ba0d68cc18406f0a562d293243c8c9;
defparam bigblock3.INIT_03 = 256'hbc28be9d78657dd1545404e625b1c70698f119ab76c8056749808cb164e1dc0c;
defparam bigblock3.INIT_04 = 256'hb2c044b0d7730bc0c5a09a08451b48292b43dcd10e45000374f6fb72f8ff59f0;
defparam bigblock3.INIT_05 = 256'hcbfb07d1755fb4284bb2db745e023bad55f3e2fdc5eb8be8d8a532a1ee68ac12;
defparam bigblock3.INIT_06 = 256'h13df86502d3fcf298c37fa1d51cfbf3e4508964570660617a1a97fef4153e459;
defparam bigblock3.INIT_07 = 256'ha6aa9c8c8cbc61a52d370f11c1265f0e173c069b36568840e3c3f86ebf445b33;
defparam bigblock3.INIT_08 = 256'h2a44d7f2b4a793e53885e1571453043a2515d8f81a24cb41aefe91602d68283f;
defparam bigblock3.INIT_09 = 256'hafc2af6fde97ad5bc353ca088b273e5efffd168b47522460c6f687bf0dcca9e1;
defparam bigblock3.INIT_0A = 256'h33049bb1d592470480f776bd1aa9912382e962eb2cbe0768c670b86017fb0000;
defparam bigblock3.INIT_0B = 256'h934d11d1279bce99140246c6a3c68983000204511fb974f790445f43cc003776;
defparam bigblock3.INIT_0C = 256'h967f8a3cc2e5b9220f1272aeba5028e58a961a86f42a27603028491110fe613a;
defparam bigblock3.INIT_0D = 256'hfb7232ff4f140665861551fc3d06287f8963c610ae96744854c532e4b9686554;
defparam bigblock3.INIT_0E = 256'h608cee249c0d7248a618df714b98454c8a0ca4bbb82b881edc694d47000374f7;
defparam bigblock3.INIT_0F = 256'h6fff1fa03bd940ef381c18d157c106d55677624be34100816098ff201246d1d5;
defparam bigblock3.INIT_10 = 256'h0162004200001160a644e68880891e9da20fd9f74aecb91b96d965f33d159f5d;
defparam bigblock3.INIT_11 = 256'hcc30a4613065050ebaa1c40b4d7014a854e1854d9791bb8c8942531491194615;
defparam bigblock3.INIT_12 = 256'h25060906cdaa94c1dc8d0352c5c65a118981875c5471677406ac80c419839da3;
defparam bigblock3.INIT_13 = 256'h8cf943d057d339974f9009ea4347cf49604c19db470ee74e2bc0e254c2a906a0;
defparam bigblock3.INIT_14 = 256'hdb849ce2604281820a20df225f550080bf7e9211139aca35efa858db6cb7ec53;
defparam bigblock3.INIT_15 = 256'h6d4168612039431062d783a8b132983a159f8133040900008109800061601b53;
defparam bigblock3.INIT_16 = 256'hdf7b6d2b7eaabb4b9e63def062f08d192eef10fbd857c9e070b7c495501daab5;
defparam bigblock3.INIT_17 = 256'hba40800274f5fb72e6ffadac6e56ad6aa8fc24f41723d767fcdcfbcaa824aed2;
defparam bigblock3.INIT_18 = 256'h8992a1a88129608aed88650a75a0c4a0276c4db5a376690ce4db902c861c5b49;
defparam bigblock3.INIT_19 = 256'he50ea252281d7fd4615f00804596ded669feeec18cfe5f9593dd3a2896db9739;
defparam bigblock3.INIT_1A = 256'h4d4240af59c412072d2545b3976a31a41e4829c000000000990837b58aa4d6ee;
defparam bigblock3.INIT_1B = 256'h6d321399b41842928916cada974840cbd44f1ddd2da9f2c89060f63d6e65116d;
defparam bigblock3.INIT_1C = 256'h3b0390ab0ac8ba197d9f9631f5bc8826d59b5db0cde4a2a054ebb637b89878c0;
defparam bigblock3.INIT_1D = 256'h7d5cf85bb217f8c96abe34408fbc936a659509c36576e73f2f8ea2353bb242c6;
defparam bigblock3.INIT_1E = 256'h7dfeb6fd718ea866318cd0a5eaa748d51bacd0f400c81800f3dfc446d5e944b3;
defparam bigblock3.INIT_1F = 256'h2447f14db95524705e8b242354204088462532804cb04e8834308f1b4d1a1736;
defparam bigblock3.INIT_20 = 256'hcb546ce124ee479d4a25036c32b32ee88a1715a228895248a4d7337aaa397a44;
defparam bigblock3.INIT_21 = 256'hf814234ddc51c760000374fbfb7053ffa0a5b2adad354da8da4606b2c72a305a;
defparam bigblock3.INIT_22 = 256'h54cdd9e53cdb5a9c6cb1412c30982e244a8555a884985b710d8543008904619b;
defparam bigblock3.INIT_23 = 256'hbb61a5718d03444ba7805821eaae4fff0000d28d6e7c0e5eda0997fcb1fde0ec;
defparam bigblock3.INIT_24 = 256'h0aec4cb3907d277aec95cecca1f5122a16c6187287c7000ac122412125db56d6;
defparam bigblock3.INIT_25 = 256'h771b064477d2e23076b2b0936f8b2c1259ce083d0b25aeac8890f6c3e9e2e73d;
defparam bigblock3.INIT_26 = 256'hdd98f43b9ecfa7312dd8aeadd6c8bcab29f5c273b2cbd7dd3dd572e407f7d907;
defparam bigblock3.INIT_27 = 256'hd2427338bd06b64cc8c0807262c8d7ffc802b72353448c2de5606bd7c4f716bc;
defparam bigblock3.INIT_28 = 256'h9a07ce4eedcd708e2531d06069f4f327813afeb0df08faf158785cc62a5cccfc;
defparam bigblock3.INIT_29 = 256'hf2e2327242ff0e9966f3774791c065af663c984bfd5ca4790d3f84d13db5971b;
defparam bigblock3.INIT_2A = 256'h015a020ab8e13e70e2cd2298ff277198f7a84428330ff32b8503b83358045dd8;
defparam bigblock3.INIT_2B = 256'h085005865b4613e11af251e946da036fff807274fffbca12e763367d6278e098;
defparam bigblock3.INIT_2C = 256'h51586f1fa91bc1207916480504b84dbe8a332509249305ade85ca5116847291f;
defparam bigblock3.INIT_2D = 256'h27d5921628e51b39999553593195adaed622d8e729b76eabef593786e5a21f1c;
defparam bigblock3.INIT_2E = 256'h23d7743f825d2ee741679e332c69b5735905e289d2f14cde48016802824c1721;
defparam bigblock3.INIT_2F = 256'h7abbb60d73b468907597fb285f14d6ec1c492c87f053e7e25e30599797ee6f8e;
defparam bigblock3.INIT_30 = 256'ha6058f3c85f3bf73100c52cf422b1277556fe8a4fd0d56c922f6e5fb851fb95d;
defparam bigblock3.INIT_31 = 256'h7742361c2b282d0e5d9386945ab822abc23b2febda84d9f846da4902c73428f0;
defparam bigblock3.INIT_32 = 256'hd07c3242b65859370e143163a25400c2000019803710d018b46d47dc412e622e;
defparam bigblock3.INIT_33 = 256'h39b0719158c91d57b195c6aac9f5cdd1089ad506cfad9dec6844a6bc0f02481d;
defparam bigblock3.INIT_34 = 256'h4ff73514cb5d16a35fccc1b5675767543390f46769315ea2f55627a933256b7f;
defparam bigblock3.INIT_35 = 256'h0cb87146f8d1084b0103db8622e31728392857dc034afd807274fffb7d5adcfe;
defparam bigblock3.INIT_36 = 256'hc752fda38cac62fa861b2ae5241c2a3070758e6599faef7614e134f68f6e40b0;
defparam bigblock3.INIT_37 = 256'h80950187600446296e5c87c5785c3803471b36cca6212ab4b691db9170364d90;
defparam bigblock3.INIT_38 = 256'h3ae3c79ffe2eb9066bc91772420b3e3d636e99a7a325699684878b752d3ea2d7;
defparam bigblock3.INIT_39 = 256'h9f629e2204ee42fa21d675c93c9d6682526fa43b1f049aa0627c95ed2ac3e685;
defparam bigblock3.INIT_3A = 256'h011f3014480098883e3acf2b865fa8577fbb249264b663504f921f565b5fdccc;
defparam bigblock3.INIT_3B = 256'hfd6fe9b21d170224d34990803b306dd4c723a10478015ff411774e832fac2b2c;
defparam bigblock3.INIT_3C = 256'h23463d43abd8c5549307c0bc365ae4f3001b4ea01a20f0473ae3b7284a7a6d21;
defparam bigblock3.INIT_3D = 256'hd5d83e3dee24dcaddb1e2df83d5dd7b7bb78adae913407e9107f90cf9d6b9440;
defparam bigblock3.INIT_3E = 256'hfffb102e25a3e60c141052da95b516dcc81d84e3209cd0a0f617b60f29d56942;
defparam bigblock3.INIT_3F = 256'he81405ade05db1726f443911740e30a2eb7a29832d20e9e844db0304fc807274;
defparam bigblock4.INIT_00 = 256'h6d7148db4002bf403a255b7b86a87e47ea99b0965bc62ee9ded2b5b767be9821;
defparam bigblock4.INIT_01 = 256'h89854a8901440000d000880b824c6b12da9022a72636a61f546e02b8964b7306;
defparam bigblock4.INIT_02 = 256'he3c941e7f14c818c9cf60bccb61e03a8e718d0c7260d5492963372820bd188fb;
defparam bigblock4.INIT_03 = 256'h0fccdca332456122bb79a6504d6587339b897deb7af224ea35bace6961ab3b75;
defparam bigblock4.INIT_04 = 256'h00010268a72fbf77bf151f48a75b27a8e3ee34e0a5a8548370e85fddf9ed614e;
defparam bigblock4.INIT_05 = 256'h1a6406e600103040a806d9a097e2cbc9bbdc4a6ca2286a8529303ae28db7c91c;
defparam bigblock4.INIT_06 = 256'hff3bf27da8b588b28666d6ebbef2d162b2d49d56e9f3fb4db3d08250e2e3375b;
defparam bigblock4.INIT_07 = 256'h696e4c8ba3b2ff53e1c3688340c9f0943ba080ccb7228a6117f3e888ee30ae86;
defparam bigblock4.INIT_08 = 256'h0395fe007074fffbdecd7ad6720040e59de28e866efaeffd6feb3fe3d7cec6f5;
defparam bigblock4.INIT_09 = 256'h4400cb0114919c268a6da06d25166cc63d27844d2465bb6a21225b18498f455b;
defparam bigblock4.INIT_0A = 256'hf937ffc3de50fc03bb332ff38364f9479190b994ab6188c644edb71e9c6d0002;
defparam bigblock4.INIT_0B = 256'h58404943213ca196b9e6624350d4406d78540ebe90013184bbd2f5207bd34d21;
defparam bigblock4.INIT_0C = 256'h74d6ffde48f55b802b6a66eb0df8df6dd48cde6eb46834a0610b78e63a20a6a7;
defparam bigblock4.INIT_0D = 256'h604958a096b7514b237eeb32f1d8153235818dead56c2824bb3ff413b0fe458d;
defparam bigblock4.INIT_0E = 256'hae1a744cff916ec3e1ac81badb7621c8fff8ffffffffffff63ff3f50dea77dd9;
defparam bigblock4.INIT_0F = 256'h5c6b585c75575e7d702202150900e041bf0583b4d8e81c1bf040380881429f1c;
defparam bigblock4.INIT_10 = 256'ha3db8c23cb0d618c72183e31606f2e996bcd725a0de408c79ab04e28d0d48e9b;
defparam bigblock4.INIT_11 = 256'hd37ab98472243797373112d94573cd08784c79626e28971d104e758f0f737a60;
defparam bigblock4.INIT_12 = 256'h701aec5a5a513834000374fcfb7231ff7bfb97f5adfddd4e1277657fadcf84bb;
defparam bigblock4.INIT_13 = 256'hfb400e1c2487a4213dca88116c18ed34ac0d07c08c3d07694c4d0c204d1ba16b;
defparam bigblock4.INIT_14 = 256'h1e1c7b05c3c68321301d7af4ec83c6e381c6e3ee8672080998c8e3e11bffd080;
defparam bigblock4.INIT_15 = 256'he5853b5956c73797196406299781f41bdc0feee93c9acf3a0000b1b640007509;
defparam bigblock4.INIT_16 = 256'hfa819ec5b8356055b2a7630ee9e5324064754a66158ce30435f81217913f8489;
defparam bigblock4.INIT_17 = 256'h2019ca33f22d53629bf768f46a5dd7269affaf4ba836a98388d9c68e723b87f3;
defparam bigblock4.INIT_18 = 256'h2bfbc1442ec6dc6d81b60800195fa8427183bc59d41960d8215858ea8e472a54;
defparam bigblock4.INIT_19 = 256'h8330cbaed1650039ce2a010881eb8fe6176eeb195bb3d8016d319b2988dea131;
defparam bigblock4.INIT_1A = 256'h390626a2106ec8bf3daecba8d8f6a85e79559a237e0f1876cffc59326c90934d;
defparam bigblock4.INIT_1B = 256'h8f3e631c7b32e7554a4c770bb6eb64baa25323b90ef58e20b78b06d71baba26e;
defparam bigblock4.INIT_1C = 256'h831a5315435b6021892c5ab93d41800374fffb72a6fffb57e02bc72a3736820b;
defparam bigblock4.INIT_1D = 256'hd36e204c93016f33d6fd63e869315e2611be148c6d58858d5748e6206f6a4d79;
defparam bigblock4.INIT_1E = 256'h850000803e2896ac9a30679613556b4c88dc8938518cfce56eaa0b296a8d36d6;
defparam bigblock4.INIT_1F = 256'hb3da38aceffaac484c81ccb90ae217d3a203366ad2a505efdc83ea480ba300ce;
defparam bigblock4.INIT_20 = 256'h4663f0216b27d8bad785580fff0d01515e9f0a35bb409467b9f09f3e954cb2ef;
defparam bigblock4.INIT_21 = 256'h0456d13541d182176f460b63ab5a045773dcdeb4ff7196de1b286737f2ccdd72;
defparam bigblock4.INIT_22 = 256'h7e336294172f87b383982bfa19538e504fffe70125ff4831501d0c8f80dba63a;
defparam bigblock4.INIT_23 = 256'h49eec74a62faf452bd31c0b5ea9491870001000400130aae332ff575caec60e2;
defparam bigblock4.INIT_24 = 256'hb3c54ccbda1ad2f989b95cc0e8247bdc38c3796d1a9043d0994fcc4d570ed806;
defparam bigblock4.INIT_25 = 256'h4bd0cc461f7c6baf99cb030bb2e1ce5785460031cea3f86a8209851736fd0544;
defparam bigblock4.INIT_26 = 256'h24a007734c59e62e9a04635b4a20881e5cd1905f800374fffb721cffb1a75167;
defparam bigblock4.INIT_27 = 256'h203cbb48ffe0800b4c693bd05cc1d9119e6169c42040899414946e68820db1a8;
defparam bigblock4.INIT_28 = 256'h0f9f963993d70e55d00047000431432eebe774530ba8e71f7cb094ef5a3d961e;
defparam bigblock4.INIT_29 = 256'h1db7d3485d5fa3b9533ebebd7d5438984d6b4f91b71731ff68f8470484f75ab8;
defparam bigblock4.INIT_2A = 256'he852a530992265e6e7d6c4a122d9d381c1634ef6be6d5c336b873b77e9466cff;
defparam bigblock4.INIT_2B = 256'hc1b0ffffffffffffffff15ff7429e4e48de1d9e91d30b1663fc1f5231ae63b84;
defparam bigblock4.INIT_2C = 256'h5d18d000ea16476294d68b7666c2267c6d22b5b6dd2a176462c1e164224bbfff;
defparam bigblock4.INIT_2D = 256'h4cb6cd8bd074153bee972bb62a68cd1eca3a9c9534ab46c294ee808400510400;
defparam bigblock4.INIT_2E = 256'hb4908c573aea9a64a54d39b98138cc3450f7362c713798d6b1df3dc6ac76f779;
defparam bigblock4.INIT_2F = 256'h6bff242551cb1379b6930eb546c77f822a916be3da1430fabfa38db9d31d8066;
defparam bigblock4.INIT_30 = 256'hed98758db1a0462c176d4d39e5226605835bf81d891cdb498345800374fffb70;
defparam bigblock4.INIT_31 = 256'he8ba1911375b0ec122b8f8b3fd9efffa4002800c935e2d8e1e958483a0051308;
defparam bigblock4.INIT_32 = 256'h0e6281786c1cc7da8b8700468000008ce400b05493fcab6ecd0a45d6511d504b;
defparam bigblock4.INIT_33 = 256'hb91f866bb2e6847b4e117893609e6989341922da809c3ce80046131728106bde;
defparam bigblock4.INIT_34 = 256'haa6d8ad8ba32d772d1ccdcbe180165d3ed4c2e0858eea2d662c6e7792b9fad70;
defparam bigblock4.INIT_35 = 256'hb6db52314680fff0ffffffff6ba7abd836a328ebf738f2214a1884f36aac194c;
defparam bigblock4.INIT_36 = 256'h1a005ff13af79e1527d8c6342bf2867968222a2f4a0c4ca34ecc528c71cf9f01;
defparam bigblock4.INIT_37 = 256'h20bb77a502367a71e5a4a80e131967fadf65b46989c628e73e251c8800006c49;
defparam bigblock4.INIT_38 = 256'ha86ba2e41c1a8145eb5f95879b388ffdb4788b6b25997e65aadd36d8f8f92ff1;
defparam bigblock4.INIT_39 = 256'h034aff807274fffb905da74de5f819f95bfeb0b9a9b9d6ffd2a0edf339559c81;
defparam bigblock4.INIT_3A = 256'h569fee3a99e1a4920d6da08a2d186d466915384d1cc55b661f031788318741db;
defparam bigblock4.INIT_3B = 256'ha06b1a2f8305dab127229f3f4faaf912d987bd9cdb6e28b8100036c221ff4d9d;
defparam bigblock4.INIT_3C = 256'h54ef019bc9e950f632d62a14f8678fc5005d440022002602c330456d0191c33c;
defparam bigblock4.INIT_3D = 256'hedbf743c5ede2bc5329ae8e9475e6f4b3ff28c6f74977b0c851117e3fddca680;
defparam bigblock4.INIT_3E = 256'h8ae85552ecbca15d7ee2ec7ebbb3e52dd9d29ae753f0365fd2bbcb7a9b234c49;
defparam bigblock4.INIT_3F = 256'h7c6d995cb24010c9ffdc15ffa01468f09052e236ce690c51afe891fba98921df;
defparam bigblock5.INIT_00 = 256'h181c0d434000284048088500fb97b0d97ad71dd11ad98fee11cec2caa4a9d682;
defparam bigblock5.INIT_01 = 256'h52cb9ed43ae9f93af69fa028ea1f908c98d1142c69153a10a4773635dc792121;
defparam bigblock5.INIT_02 = 256'h8cf420167499bf4d5838dad41f7a0a74995245fdd623bb9b40ab9e330ad7d769;
defparam bigblock5.INIT_03 = 256'h2f885126415b0354ff807274fffbb9f11c88bf741f5cc84a8d654908e5594e9b;
defparam bigblock5.INIT_04 = 256'hed613bd015fc5ddaeb6c89d8a8920ded288f1cbe6ce62cd1724c18465b6a2663;
defparam bigblock5.INIT_05 = 256'h0a3e3a3d4b67315f20d95f5380921d5034506835f629ee407ba76db7906300de;
defparam bigblock5.INIT_06 = 256'h1d28262d35830d2928178aa1040da51b9ce85100000164120008abc04f50137e;
defparam bigblock5.INIT_07 = 256'hcf4b482057c61c23d4c89a7de2b949978c6c06a3cd67823b1bd1eae4265085b4;
defparam bigblock5.INIT_08 = 256'hc0a7b8db855f737a9042eb14ca2e22b952387bfb5b9d3503e3d507982b05bc93;
defparam bigblock5.INIT_09 = 256'h189a194dbf8b6db682630000fffcffffffffffff7fff2ccdad6a6eaf1b49ac73;
defparam bigblock5.INIT_0A = 256'h8000580000003d337330561b729d963e80bfb4a25c93b2ce779f692084eac3b0;
defparam bigblock5.INIT_0B = 256'h06361146ffa3db841955698d241616363e490dcaab525d636a58daa0c8c21b18;
defparam bigblock5.INIT_0C = 256'h0885e873f84652b15b43349e881d525acf66ae88a9cea6edcf44a127b766c432;
defparam bigblock5.INIT_0D = 256'h24266b6923a3147861ec49db0344ff807274fffba185a8b4a430cec74c700c44;
defparam bigblock5.INIT_0E = 256'h00805a68fd9d7a5d334bd8f4557efeca1ec1a8918d6d209a205e6da6c919720c;
defparam bigblock5.INIT_0F = 256'ha00630a4056796ba7f66a0cdd9283c4ee597283a66bd13ed4f0eae1f36017fff;
defparam bigblock5.INIT_10 = 256'h62803bcf6760da54e91ec8d5830825de016ab53a1418520d1e1847512f86211c;
defparam bigblock5.INIT_11 = 256'h6fea4039a9e7636d07c8e4c1d758d510dfe20162decb297e21120d3d98e5fce5;
defparam bigblock5.INIT_12 = 256'hfffffffffffffffffd3f7aff5b3b886adab7c83d1b97ecae1667b4a4393b6214;
defparam bigblock5.INIT_13 = 256'hcda4a9e8a09e0ab4ed5be5f199cc50b5dbef8542a85b6063db6f4eb62000ffc1;
defparam bigblock5.INIT_14 = 256'h47f562f729a162ff6ab9e99a2359758bf4f1478000053050ae948820338070e3;
defparam bigblock5.INIT_15 = 256'h10c53bbb305abedaabac0ea27d27f769733a247af185a256fbb2fe709331a544;
defparam bigblock5.INIT_16 = 256'hfe65b862df75d58abf9b88dcddba9cc7c674574664a9c832a22d7d00be98a9dc;
defparam bigblock5.INIT_17 = 256'h6d46f507940b24697b6a26a31638512b415b036efe007074fffba03c60af7934;
defparam bigblock5.INIT_18 = 256'ha43907593a04f746fffd02044842c7a7cbf09ee5416994b198340d6da07824b1;
defparam bigblock5.INIT_19 = 256'hd6b8333f07aea00002042aca95d420cc0c20ab1f13a0ebf7bbecb03e504e79d4;
defparam bigblock5.INIT_1A = 256'h5461cd8ac136b38410d5cbb39fc8ae9326b24cefed2c84a1c956bd3a7692693e;
defparam bigblock5.INIT_1B = 256'hb4a1ccd3bc9222f6044ea8131c6955aa6d8296c25aed714261fbc4813e2728e5;
defparam bigblock5.INIT_1C = 256'hc50cf2616ef9e126a4df7a0cd6bfb6614f8fb9b40fedd6bc0bac3f7f57f33d54;
defparam bigblock5.INIT_1D = 256'h09a811523bb889b4152bafa06946371b0021577f07145be1a8e124d18bb136c2;
defparam bigblock5.INIT_1E = 256'h8a89bdace120e9c326dc00c71218848057487ec37f88f0ecd9c0ec36ea11e8e2;
defparam bigblock5.INIT_1F = 256'h0361d4c4e8756647c2325432ab29717ab194e9af0bbae2e3ffa1bc93052d5fac;
defparam bigblock5.INIT_20 = 256'hadff15c39b0651f7bf2a4370feb2d9cd75c74213fad8ffac2f60d37a482affea;
defparam bigblock5.INIT_21 = 256'h6da48d8d5ae0e62c156c0cf1094c6a15e37bc8252b2d5b312a41800374fffb72;
defparam bigblock5.INIT_22 = 256'hf290aa6ae46d189453011a81ae71e3ce12a256d109f04081e2c42c1e88c3611e;
defparam bigblock5.INIT_23 = 256'h5e8e38230640a00080a414e9ad74b333465cd907747c27c9d3948dfa91a2c242;
defparam bigblock5.INIT_24 = 256'hde3e7cd3841645ad939f352910db3bca115673f356e795a90be99a56a8744553;
defparam bigblock5.INIT_25 = 256'h0639aa9098faf88b4b50cc1b6c8d07e76cca6b7cf80efeb00c172711de3e7299;
defparam bigblock5.INIT_26 = 256'h5fc0f6a18c70021545c3d55b0233a1685b8a127d72e8a9c72d37d5aaca2bdd2e;
defparam bigblock5.INIT_27 = 256'h654cf0ed4389457fca3ffc0f225805d04ee639f09bcde265660757a238db104e;
defparam bigblock5.INIT_28 = 256'h8ca960b1298ed1560f37c3b9cc54b5a75c1a23cc0b681ba802dd300000251478;
defparam bigblock5.INIT_29 = 256'h067e28c4e55b588a5fe894cf7b15905d11e5611ebd08559e26e2ad80f6697b4c;
defparam bigblock5.INIT_2A = 256'h800374fffb72bbfffe55165398dad2ad6b98a18890743b63f1c71746ce0df911;
defparam bigblock5.INIT_2B = 256'h8b7238d113086ddc7a8d1460262de16f0c6846767720237bf822884ddbb9c060;
defparam bigblock5.INIT_2C = 256'h39df2f7adec5e69988855187e5a557a6e38d2d2824000e48d887e15abbfce774;
defparam bigblock5.INIT_2D = 256'h734cb2ad3c35bdba4602000004109490c4658711d5b8d8d32db0d81dff2528a4;
defparam bigblock5.INIT_2E = 256'hbcbf96e19ebe9453449957144b50f1b792573462183e72ea5ee46d8363d64271;
defparam bigblock5.INIT_2F = 256'hbdfd3a9aded572cab4e3caadfe5e65e71b88fa15b24db49776a6d0607d7f1a47;
defparam bigblock5.INIT_30 = 256'h52c80a2f6590a3cae46d1024c76e7aed3a1bf5fbb8d30a2d9fff53e63d91c28b;
defparam bigblock5.INIT_31 = 256'ha3b397c4000285a048028217c5f8bc14a5d858bee21713ca5d4ab46528733991;
defparam bigblock5.INIT_32 = 256'h6a7b75d1b4a975a583cddad31377ef8b54d96447066b87bb2ba5d37ac158224d;
defparam bigblock5.INIT_33 = 256'hbd3198bf1f1c0cc1ef18b62800e4d07c6ebbe68232785819a3e94614d67d73b1;
defparam bigblock5.INIT_34 = 256'heb2c5b394a49800374fcfb721dffe9ebf30ed6d924f863017a43d8abd1f06261;
defparam bigblock5.INIT_35 = 256'h52461623abd4d0e5a9db93096da8998defe047a4136d0ca12326670d636b7821;
defparam bigblock5.INIT_36 = 256'h9b0a008a16355fb12a01f2a130a3efae4f4d1e13f44ead625247c2cbe1dddb9c;
defparam bigblock5.INIT_37 = 256'h214a57b64912c595b05a7d35613c5b980b15784f0d61f4e9073142209b2cd077;
defparam bigblock5.INIT_38 = 256'h06e5803c56c988267826c75450faf95bc38e5d503c64efb09b88ae5857954d5a;
defparam bigblock5.INIT_39 = 256'h50066f9f47df650f0ad557731993d2b64ea9cdfa952330f1de6d2d4788f2675b;
defparam bigblock5.INIT_3A = 256'h196560899c8077b46db8832420004f0828bfbfdb676512b5073748e923e53fdb;
defparam bigblock5.INIT_3B = 256'h049c00405e08d1a5aa17c872b63205588172b93a1f21ada87cd43c26d6884e49;
defparam bigblock5.INIT_3C = 256'h641ee0c39de3af2c0950658dc5970d3b2884076e37ac291f194c7370c65a9252;
defparam bigblock5.INIT_3D = 256'h52ddda1f32ca2a4d72752ea29ed51111f6ab141159908e1799331858535910b1;
defparam bigblock5.INIT_3E = 256'h570042bbc822e95bdad11b44800374fcfb7032ffe5fce3df3f6db6cf5e6b115c;
defparam bigblock5.INIT_3F = 256'h5c6d71b7012400006b08e8f41d7ff8fdb4a06d5c9c8cbae04620136b4c49c70e;
defparam bigblock6.INIT_00 = 256'h00a179579a672a3a3c8b064989c3b566b2c8ec4ad1c948466d544176451ad07d;
defparam bigblock6.INIT_01 = 256'hb0b70913545078b91a903d78b22a97c1a40d79a25dd8c3028b2aa609a474000f;
defparam bigblock6.INIT_02 = 256'hff6e3d2896cd1f9dcf843b6743fd51a96ad3d841393b3d39d3f9c9d1dc650633;
defparam bigblock6.INIT_03 = 256'hf6c16044c94fefa11d8a1c728d55cdc8cd4d302ae9979249f67745a2ba06436a;
defparam bigblock6.INIT_04 = 256'h0a85dcacf1ea3dc63abdb0483576a492a000fffcffffffffd7ff4725cdfff7e0;
defparam bigblock6.INIT_05 = 256'h46e8de4c1b9b9b5b0123704083408d1650c6ee269dca02a707f287ba8c5920f8;
defparam bigblock6.INIT_06 = 256'hadf65ded6683910567e5f987206f0cb13bc590e6e5dcdd17697693fda4d0e174;
defparam bigblock6.INIT_07 = 256'hfbdd3810c865ea54952c0b3003e5b5fe4e8beef9a228f6f2c3ff79c0494b7bd3;
defparam bigblock6.INIT_08 = 256'h66e70905820b25077b3a29c31d68b1eb45590370ff807274fffb7ca3d35a224f;
defparam bigblock6.INIT_09 = 256'h1d1e07d03cc4e743238d2019e900352cfed6d9db75ab1c38e8060dec809cb0e7;
defparam bigblock6.INIT_0A = 256'h2a0712e91283000055003ae377540082f6cd1416836f62b6f8d3b0865b3a73d7;
defparam bigblock6.INIT_0B = 256'h347d1a5d333249149d3b3a58abafa7093d98ddb22e9c2a58771d11ebd9fac392;
defparam bigblock6.INIT_0C = 256'h1fc5dc3042e0d8296b32c54592e919861501f6f033f3bd59c5eecb58a94b3773;
defparam bigblock6.INIT_0D = 256'hbfff55aaddfd0d338df77ec009eebee61d90f71f5ca2bcd4683cfbdc036a7dc2;
defparam bigblock6.INIT_0E = 256'hc748477fff49e70a0da5bfea37388eda116d384aa0737241c6ca5491fff0ffff;
defparam bigblock6.INIT_0F = 256'h0ec1ce84a95237098ba382dd7155c782580f9707d01d0003b800c61e592e34ee;
defparam bigblock6.INIT_10 = 256'h92580619ca8b1dd721c834696981a67829eec54ce40496954860c9bcd1e63c70;
defparam bigblock6.INIT_11 = 256'hd002483d1ad8b68f0c34967926181735ec726579ff32c7192c919116116b3bbb;
defparam bigblock6.INIT_12 = 256'h0d6c4090a4b366e77d03284b0d855b3725631798b1884d59037eff007274fffb;
defparam bigblock6.INIT_13 = 256'hf51ea8e88421964aadc9ad0a1feec7a0c3259492f230b38ed3d658680969dc93;
defparam bigblock6.INIT_14 = 256'h99b2a562c440ab84721e57250000e500fc1c5cc485a64f9f2f18d51842e64385;
defparam bigblock6.INIT_15 = 256'h7d195b265ea59fdc9018adfd5b48168412ef1d225160066a96c63dbd95720e8e;
defparam bigblock6.INIT_16 = 256'h83246103dec09e45013e83413e8d67309950d5228eb33219e2fc4c5e7103bc82;
defparam bigblock6.INIT_17 = 256'ha6da0bfff8405fffcf434d3a5a1733c3e921545ca93d237381ba2f7c63dd0569;
defparam bigblock6.INIT_18 = 256'h412038680e65b81a48527b5bd8964e1b1deeda43810d0485212c0aa4f10e0924;
defparam bigblock6.INIT_19 = 256'h75ca3b6b4a8bce0f8ec2c762750c0aacae154e5660f3c3c5426124032aad0000;
defparam bigblock6.INIT_1A = 256'h50ae976305cc4d99fe1a39206f7609cbb9f7fa202f97136f9c4e8286e4b5a58e;
defparam bigblock6.INIT_1B = 256'hff807274fffb34cdd42eb0e26182801092119d0024efb61e58972f763235b4b4;
defparam bigblock6.INIT_1C = 256'h3ccb8ca1c8340d6c607d20756666e4e3064c05063b3323231f98998845590364;
defparam bigblock6.INIT_1D = 256'hf35e124ba345e27131abea472e4c1a038b9cb3ccb612fdd1c105baa05a93350c;
defparam bigblock6.INIT_1E = 256'hc75a3b1538d9adadce66cca4b76b1b4a2b4200000060cc0a333f34a935bf687c;
defparam bigblock6.INIT_1F = 256'hbd965b5d408713428cd51b54c86edb84c7954eb85cdbb9a39ead1c3a09dc9ea8;
defparam bigblock6.INIT_20 = 256'hbd5b10bde77b79430bf835ad2799c7b13339087a8ab8534033bf9e322efe3fe5;
defparam bigblock6.INIT_21 = 256'hfffeffffffffffffffff5257266032029d2cd8298b4a3a69901ebe6a14b2dfcd;
defparam bigblock6.INIT_22 = 256'h0ee58b60002a6000d20473d4d73841d117db4b8cb6014446a89a1da8bc98ebee;
defparam bigblock6.INIT_23 = 256'h49665cf27138f232d6a2792186c8c0de02b16b1d25e6db9abd6fca738e712a79;
defparam bigblock6.INIT_24 = 256'h7b77df585b3b6ea3b4fca3133e89536d28d71ccc2c3189dd13dce289cbacbc42;
defparam bigblock6.INIT_25 = 256'h99e93d58034dff807074fffbf7c3f23e7e79bdffa57efc7d1ddf29ff67cf72fd;
defparam bigblock6.INIT_26 = 256'h80683d8960f0a740986158640a6ce0921876626644e3580c2cc27b1624c31bf8;
defparam bigblock6.INIT_27 = 256'hf035db04af5ed87f96fad0f9ebc1be6aaaab25ea16ca7d41f0343ff023ee8c59;
defparam bigblock6.INIT_28 = 256'ha905c998ac6c9104819349d04152dccda93338049a5083c9005200002cad7e05;
defparam bigblock6.INIT_29 = 256'ha25e0d4b258ea865bd474eb1863863a6a09188921703e10fa26e0a84e47a844a;
defparam bigblock6.INIT_2A = 256'hec87cf15b3e8c1645eb66a99e1a71990927520af5ab6772319640ccf140c75aa;
defparam bigblock6.INIT_2B = 256'hdfe78d6a4ff78fbf47ffd69f8861dc55345e9a1da56756efeea2891d4cd3e32a;
defparam bigblock6.INIT_2C = 256'hfffff03f18a3f838fd40d4fe29554819ba085ae4410a051b325ad072e719aa14;
defparam bigblock6.INIT_2D = 256'h45a300fb010d6698fce042489f0e423474a44d857a14892990910e6a2c4eff67;
defparam bigblock6.INIT_2E = 256'hf354a1aac5717ad87a3ac7e55abe677648660e0f7df6b094139769961368b2ea;
defparam bigblock6.INIT_2F = 256'h121941fb2817e61e58b9ae4b800374fffb72b7ff0883da169026705a393280e2;
defparam bigblock6.INIT_30 = 256'hc98034b4a2e7be801f466b4b2c0a00c69860ec4a5d078020f4f40d620e39e920;
defparam bigblock6.INIT_31 = 256'h5d9c293429d61d67b0adfc9f154509ee8e98902e03a10fd67b538729872e11e0;
defparam bigblock6.INIT_32 = 256'h58fd212800c909b54609f1688bf3485c470575bdcb0a6f333fa4168d887aaf53;
defparam bigblock6.INIT_33 = 256'h9f371a8c574e86ab7a28a6d555cb4356b98c8a407834a449741010c2624598c0;
defparam bigblock6.INIT_34 = 256'habd265b672925ea5131d84478fc988c9f61a4edc8245132b538ed0cfb11b8384;
defparam bigblock6.INIT_35 = 256'h0b9fb70e7cf1d7a3bcec235a7543642ec8e5c6c11adf9ad97546dd3cda18bed7;
defparam bigblock6.INIT_36 = 256'h4359fec2ffffe07f0c176eea21ca3063ec2ce7ffccbe76e60fa696d7f9d864ff;
defparam bigblock6.INIT_37 = 256'h13b439ce58911a5552e75d224d56d65ca5c10e486ccb46905cd0550aab228f47;
defparam bigblock6.INIT_38 = 256'hd4750014ee567ea6bd0e7c58d4db550d00f2cc23595b2a9f472b7bbe23c8fc42;
defparam bigblock6.INIT_39 = 256'h915a1abdb000d2c703ca004261e05696c43f800474fffb72b4ffa6105c07dd8b;
defparam bigblock6.INIT_3A = 256'h15524e72a1001160894e684c974638ebab5c7cc500f31ef02b4b0e8f800119a7;
defparam bigblock6.INIT_3B = 256'hf3d53a3b207ba91a6beeffe1dcf9e16a8ec5683ebb7b97a9aa5708cd758d212b;
defparam bigblock6.INIT_3C = 256'h39cff7dcb7a4394f7becdf3e13b5a99f801cab765414f1f25f2d36cdc543d455;
defparam bigblock6.INIT_3D = 256'hf30a10094744cb765dd8579452b91a0eefed7f95b6db1a8d0138400116c1ea83;
defparam bigblock6.INIT_3E = 256'h48653913cac38c413a850ae70c40955a4e97226636f5b205493414bd62ec4b59;
defparam bigblock6.INIT_3F = 256'hc9ed3189436bf3ae237dd82893820ed84c9df6120e360172fd31bcbfbeb25f0b;
defparam bigblock7.INIT_00 = 256'h50bfa06d61cedd95db5372a3acc54815de7a9455ef212c6534653bddecd3231a;
defparam bigblock7.INIT_01 = 256'he3444672c7ddcab29cc9daaef576a349bac1264d34bfe36dd904740657eb5bfd;
defparam bigblock7.INIT_02 = 256'h2914f88bd4b88a49419351c48c2257564e38fa6f93726c4797a64824eeeb252e;
defparam bigblock7.INIT_03 = 256'h690d4bc8a3244b794c2d9400cde2e2fb0a1e3100de67243c80037490fb72c1ff;
defparam bigblock7.INIT_04 = 256'hfba5747f2afe8fd8e08916657a5d987ba3ac18731ab7f8914b23a8941119ef28;
defparam bigblock7.INIT_05 = 256'hc66f3c5e906f54dce1acdbabca6e7cf7476dce27e34959c7c762c3f9a59ff447;
defparam bigblock7.INIT_06 = 256'h5d50d147a7d3abbfb55a16629c042bf8b692d3cd4356800371cdfdd0bd1492bf;
defparam bigblock7.INIT_07 = 256'haaea77d6a46f100b9e54cec7447c32ba5a53038792e8d883e44f6646e47d8ac4;
defparam bigblock7.INIT_08 = 256'hd11e32eda4bb4da23d7f6fdd87508ee6a0d8558881e31116eb1865fbc4c9fb04;
defparam bigblock7.INIT_09 = 256'h75552dc2f13affad6a7954dc9137b0987cc5ecd6b2a97d1aa6652dde90f486ba;
defparam bigblock7.INIT_0A = 256'h4c894b098837f848ba198c0cbac555ec1a94a9d74917e6dbac5a20b445002e85;
defparam bigblock7.INIT_0B = 256'ha8ae266153c66f6a3a5623b9fc0d35772f0f4219a0cfc79009a20027b700526d;
defparam bigblock7.INIT_0C = 256'h749cfb70cbff354ae58bea0f81365d54fc390e4814fb7bb5b444b19e7d29e87b;
defparam bigblock7.INIT_0D = 256'h60480088efb46b0d5408a5bc277d0bf52732ed00837bda1be91b5f69293d0003;
defparam bigblock7.INIT_0E = 256'h2b594b8f6acb1fec41c21496f075a4ecbbbd4e7c7ef25afc641fa6d41d5ebffd;
defparam bigblock7.INIT_0F = 256'h4e81a1930afe396354ec0ab478c1cf7a08a8494ad3f46da5c91b158121e29d91;
defparam bigblock7.INIT_10 = 256'h0e08bce20f5d476c79d1267a63fac8bfbc8fe5ea0da1a82040204e3604c94b64;
defparam bigblock7.INIT_11 = 256'h353a675aa36f78154478d83add1f30a757d84c3f8aea6b71a246d7afbfc72d1b;
defparam bigblock7.INIT_12 = 256'h0965cc43810bbbaf4b42fecfcecc992e2621e7d19bd01915209d377ddff83b11;
defparam bigblock7.INIT_13 = 256'hd908e2690022930a86acbd5d2032b4f849d2c89c6cfd38364bb9b6db0f314019;
defparam bigblock7.INIT_14 = 256'h4ca9d7f85acb8078224bc5b3d433eb5faaa7099594530d8091b894eda9b4053b;
defparam bigblock7.INIT_15 = 256'hb9276dd06795fd89743727597d34374007d1eafab2903f8a792ff99f93873309;
defparam bigblock7.INIT_16 = 256'he9892edd030ba9007274fffbed6f57dff3e62c76453696efa51d53f7c8a514be;
defparam bigblock7.INIT_17 = 256'hcf004b9d9b606e8709c0e8200deea867945877a4e957340b04657bba1da32d9a;
defparam bigblock7.INIT_18 = 256'h9469c79491e0c20d77d557d0e0c62d4a22769b68535bb06eb4ee1b6d09470751;
defparam bigblock7.INIT_19 = 256'h9cf98e439755c3d21c972d3b2a45c2b238f427bae7ad2b97dad99d6580043916;
defparam bigblock7.INIT_1A = 256'hbca913beed12afe536abb66198870856757ece94260c75f32827c895b514f4a4;
defparam bigblock7.INIT_1B = 256'h9d281cd915a177ba7f1322b7723ca683c31c5d21ca137f4cb9554cfc4ff9c304;
defparam bigblock7.INIT_1C = 256'h044b4748fb7d03820ebbbbd4cf57e964ee289703662701536d2cd91b4a856124;
defparam bigblock7.INIT_1D = 256'h2c75b91871e6f29f96bb94fa071dfe8fdbb65fb8495fa0b74358288840008512;
defparam bigblock7.INIT_1E = 256'heaccd43d19fe6d992318568a038b5756c50287cd43312b71756e3805f9883814;
defparam bigblock7.INIT_1F = 256'h4e46a611008928f0b03524f9d86f5ac60b920bbde516d2e57746cff9e9e8decb;
defparam bigblock7.INIT_20 = 256'h7bcd1e232afa68cc4d5e0308b8007274fffb55cae85f08c56b0471183ce2db51;
defparam bigblock7.INIT_21 = 256'h954254baf3c648e08ffbb7d1de918e1834128defa875087a79a6512f020c0022;
defparam bigblock7.INIT_22 = 256'hadcf2c90040853317dc35247b66d47342e7b7b94acc66ca732bed1b646890025;
defparam bigblock7.INIT_23 = 256'hac588a234655e22eee9ba09747735343a4610c7ae5ea9a28345df1e9145ce5ab;
defparam bigblock7.INIT_24 = 256'h969036d7d99231220022e04cd274e1775352c8bfa2c2ef1ea09af96dace8046c;
defparam bigblock7.INIT_25 = 256'hba844008adb410e3892082b11ab5f1c4e9ac7ee5db12c72186f00103613da149;
defparam bigblock7.INIT_26 = 256'hc3068acae0c50afa1c018f6deb5de5faa4b8b40cc5c76d29cea56f7d16554cd5;
defparam bigblock7.INIT_27 = 256'he09ff5af19c8bd969105c5b32b34a79788c7f19a71fc07eea1c00eeff88de960;
defparam bigblock7.INIT_28 = 256'h159babd691b494dc9c2d40066e3b9fd89de1bf7a87eaeadb40d205f8ee76eb6b;
defparam bigblock7.INIT_29 = 256'h0e1b84e1002692244f48c60bc7065c63e3f8465cfe18e83a706e3d3e8c9257d7;
defparam bigblock7.INIT_2A = 256'h38df020b00237b9d1e833d38e9e541dc02e4c3807274fffbe4d6563ed6226c9b;
defparam bigblock7.INIT_2B = 256'h684d4b3aa28cbb5a6ce4a4931a24211b50d3cd9109a074530c6e6085acb67344;
defparam bigblock7.INIT_2C = 256'h7d9b3fc6727a97fc11d265cbe40b50d60fb63302931b62a8218fd9da543ee55c;
defparam bigblock7.INIT_2D = 256'h6b5948db1a6528bbe208154d76c613a8f04f9f0eceba7418caf6e84d6fdcf3fe;
defparam bigblock7.INIT_2E = 256'hd1ac0005c022505d2e1bb07cccfca31fa0b6f21ce906b210b711080c52ebacac;
defparam bigblock7.INIT_2F = 256'h4ca70a6cde388407125c181d0c7f334a54475d614c9359da7b16667b54b91ba1;
defparam bigblock7.INIT_30 = 256'hee93dd947f9c4a4caa8b5a8c7a6a9e2a744bea3502ebddc4a15daefcaea011ca;
defparam bigblock7.INIT_31 = 256'ha36d9032e008d9bb6fb8fe79f12039334366dd0d5350a221e8b735ec771fc81c;
defparam bigblock7.INIT_32 = 256'h20805f401600b6ee964379ba10a2382089401706456298ce4c0f027fe67db4dc;
defparam bigblock7.INIT_33 = 256'hc5bd990f31efbb8ddd782da015323cdf88d675ffdd81bee10b3fd4affbcc0aa0;
defparam bigblock7.INIT_34 = 256'h2884a4af75a7d93d1e4b00c5bbad1fc2126a692c49dd02ebd3807274fffb3839;
defparam bigblock7.INIT_35 = 256'h92d9d35cafe5179a1e116a1f63397f73a244c4e43abe2539ae970990b4738dee;
defparam bigblock7.INIT_36 = 256'hcb76184b037e87e343bf27f57879a1baf5d29f4ee5e54cab893be3fa65b3d232;
defparam bigblock7.INIT_37 = 256'h457584d600000024ea00449f83afe6d40758f5708e0947ee2492538922244001;
defparam bigblock7.INIT_38 = 256'he2a29a46459bcaa941c6496407032b97a2a19835b8b97c7eaf50ac6c652789e3;
defparam bigblock7.INIT_39 = 256'h2a397b8f6fad51dc20e4f5e6dfb5b79aa76908a8c7e2ac66cf765a850eeff4c4;
defparam bigblock7.INIT_3A = 256'hbb96f47797d30d980d8db5afb1b157e2ef6b824fd9ce97d65769f7dc6792b3e3;
defparam bigblock7.INIT_3B = 256'h0091a5801f9004c1d0f41c3549c5ca8120c46a772492405106f8b149d5fbf45f;
defparam bigblock7.INIT_3C = 256'h697e45558abd54bcb6ef35bf79fc1442203db1ebe8565c85180b8063202c0000;
defparam bigblock7.INIT_3D = 256'h7074fffb4af54aa26d771bc11d3f5c46f47cc1f2590944dd7eefefc01388cdf0;
defparam bigblock7.INIT_3E = 256'h9879f411076de85a20726f46353b0a0c00c27b7a20833c5ad1854bdb0313e000;
defparam bigblock7.INIT_3F = 256'h2100ed05e66aeb22a7978184c06879b191799f91e267d5cdacf649bb72b9b78a;
defparam bigblock8.INIT_00 = 256'h7de83a5f3ba1735d0572cc4dca3b1581d5f5040f580060554c79c55d1380e466;
defparam bigblock8.INIT_01 = 256'hef8c22345ee95a32cd4261f435bb5a39f1daf7be942eee9074dc00060800453a;
defparam bigblock8.INIT_02 = 256'h331cf2762dcd31f23f0c32b78c67d57684a8bd3112079ce442446ff4c322b644;
defparam bigblock8.INIT_03 = 256'hb223867b244dde2d82e53e51986d401600d4edc56d0de4bcf8df864b78f0ff99;
defparam bigblock8.INIT_04 = 256'hb02b339e3e8405cf4ec6945a567bdfddffffffff368deddcd2fff4775edd9fab;
defparam bigblock8.INIT_05 = 256'hbbe2e1431beb1f54faf422605632b9200cc1a5f10b8a0d2d0000f68062c3422b;
defparam bigblock8.INIT_06 = 256'h136aa80d0216385ff8280963907e16eb69c2ee421f3a265653d8a05c500e0867;
defparam bigblock8.INIT_07 = 256'hd949854e000374edfb72a5ffcf3223531ebde67b18a61eecccbd411cdc540330;
defparam bigblock8.INIT_08 = 256'h5329aec30dff700a3324aca45d877720262033654d2d46482718a1cb4a15e933;
defparam bigblock8.INIT_09 = 256'h753ac1c6558a108b1f763fd5d34a51b6512805ab2a9865d1f4ff4cede211fc0d;
defparam bigblock8.INIT_0A = 256'h08a75d468ac9a68451fbb39e4ccf386da0532e2ae95600300000589c26092505;
defparam bigblock8.INIT_0B = 256'hcfddacd165e5c46d1fbfacfda376bbcb2a01befe3647b16a004a5b59ca716cc6;
defparam bigblock8.INIT_0C = 256'hfff3b55f24dfdef3fe6228dc997fbe67bebe5944ff1578313cf0a7f95dbbfc83;
defparam bigblock8.INIT_0D = 256'h8206ffff038454abd6bfe4eb11ff4563242d1d2d2e73fcabfb4f77c717a7bbe6;
defparam bigblock8.INIT_0E = 256'h4d6218d60000010007b4f7619038536b2694a3f24c7e6342d0051059b4a7e24d;
defparam bigblock8.INIT_0F = 256'hfe00d9d8724af227025ba9bdd6b4309f3e9723c327159f0c3ce39cc09f36a2a1;
defparam bigblock8.INIT_10 = 256'h12a2d88eca10bbb98ade7ce23cded69d2c66b54b0fb8c52f9330dfad9b467cbd;
defparam bigblock8.INIT_11 = 256'h21db5a15e933d8b17134800374f4fb72acff973f7befd14a0d4fa5a3ed721425;
defparam bigblock8.INIT_12 = 256'hfd418d62baed55e0e64ed47f295c260cec4c57066d2866240d624cd926601224;
defparam bigblock8.INIT_13 = 256'h264120f1b66b36b5ce2c42fa3b683a1699ea3460dac8693464638346b325c182;
defparam bigblock8.INIT_14 = 256'ha4ab8c02ad9ccf581d4965195fadbb3e3b2dec6b47a98474f340a82f00500000;
defparam bigblock8.INIT_15 = 256'h76179eca1d6df64adccbb64effb78e8baca54de94b6aa3e73da4e4076ecb2b4f;
defparam bigblock8.INIT_16 = 256'hfd6f141be7c6e7dee7e998ebd1488b512b99e52618b106350dc375a478e0552b;
defparam bigblock8.INIT_17 = 256'hc7a79859d1962d24fedcffff55ff49ddd5cbc32bff1e0db439ac0cbebcf5afc0;
defparam bigblock8.INIT_18 = 256'hcb4201649e9a5ee07a7d1fa500060000106bc595bf4f06ad0fd4914a93796aa5;
defparam bigblock8.INIT_19 = 256'h138ff573611c9e80d61d33868c2a66b29c755e12480c86b3e8a02351c8e74ccc;
defparam bigblock8.INIT_1A = 256'hb4474a21ec99079a3e9dd073a665129ad1711765dfc96e0f9c95d2ae60772a63;
defparam bigblock8.INIT_1B = 256'h0d718634f719a1ea4a19ec34d799c14c800374fffb727cffbb1e9d63998bc72c;
defparam bigblock8.INIT_1C = 256'h7d296e8f2a71ae144744d62841e44548f168e1b766186bcc63076fe0e7b0275e;
defparam bigblock8.INIT_1D = 256'hf48255f10000e700a2946e52834e936258901c8bfa94a336fe2bcbc25636d757;
defparam bigblock8.INIT_1E = 256'h4f96a4aec4c6bb7a33577b10a2f25fc3ae38c71e547b886c813ea78c1ef17470;
defparam bigblock8.INIT_1F = 256'h1826db3c41e519b0ae82d2d4bcbfc42eb4a5c76ad670cf651233618749fb5b3d;
defparam bigblock8.INIT_20 = 256'hb1fa20084741b2493fcb98a4357b3223dd2dbc8e10904e392745b9c11ac65cc5;
defparam bigblock8.INIT_21 = 256'he303152c88e0e0eb1891921c8c90fa8cfaafffffffffbfffa4069ef740c56ce7;
defparam bigblock8.INIT_22 = 256'h313a710d8b483561461678a972714de68edaa0e902b2000026201fb84ca52d71;
defparam bigblock8.INIT_23 = 256'h15b14c7d309231c48504b06914473c5abc535e42715499425613c22ce2218045;
defparam bigblock8.INIT_24 = 256'h15f1e3290a993fabe5e794c5d9353a4cd252d8d0e56c5e116b77b5398accf3cb;
defparam bigblock8.INIT_25 = 256'h752067a40b5c4d798918e31981dafa19ec1b5719b74d800374fffb701aff142e;
defparam bigblock8.INIT_26 = 256'h888d8607bbf9866ef30a08567195b9ac8924216e39f2bd51094097a56b886387;
defparam bigblock8.INIT_27 = 256'h44da816e6609da1c7b0700014300988db9e7e0a915f015939e8df38aa0a81d3a;
defparam bigblock8.INIT_28 = 256'h77c73e1b3b424089636c478535051813d9965f745d80230c1a347cc7f4c031fc;
defparam bigblock8.INIT_29 = 256'h70352f4452351909625530004a4457331027bdbb911f0ca8f0999c9a8ea208d8;
defparam bigblock8.INIT_2A = 256'hdfffceb8508a8d25f3f7ff67ea95cfdfda7485e171450bce397f6b329f84626e;
defparam bigblock8.INIT_2B = 256'h41e7ac7a3438e4dd7201f9885a21cd606104c0297f05ffd5ffffffffffffffff;
defparam bigblock8.INIT_2C = 256'he9a5d488e01abb8fa350ed91729fcd366391aed58c9551a2752905b20000e440;
defparam bigblock8.INIT_2D = 256'haf93c73636312263115ea65c10486b4f8224fa4a719bd58b911c09f0c48d018d;
defparam bigblock8.INIT_2E = 256'h7274fffb9679d7ea56885cdd132dcfacef657d58ba5e31e8b22748d023893883;
defparam bigblock8.INIT_2F = 256'h18a14896076be067a46f5a67ad07504d2589cad219611e9899e649d603acff80;
defparam bigblock8.INIT_30 = 256'h1a88831be5e7f66c2526eae402fe40006c7af1e5e871e218bbeb66f49f46395d;
defparam bigblock8.INIT_31 = 256'hafe834e7119ad826ebaebf1e1559e2b10075d20034aab8347a59191f3cca8b30;
defparam bigblock8.INIT_32 = 256'h18be897109a850f365d23f87607e95fd5f2bb89eac3b88b2864fd273e366aa8e;
defparam bigblock8.INIT_33 = 256'hc53e92ac96b29c72ebcf26fb54bd3ac87158ebfcbf6c24586593b8f16870fab1;
defparam bigblock8.INIT_34 = 256'h4a3b576d1d48f2bafa1e9ae3c549af31ece5c9dbada275bf325bbf4d7ad5fb4a;
defparam bigblock8.INIT_35 = 256'hf464ea1ab03cc6ba58dd58b8884aae9d7feafde3ae3f5bd7e9eff623de3b07d7;
defparam bigblock8.INIT_36 = 256'h25378e4d09969035c62d28c914680038000062600a457199c6f3838ef37e01d8;
defparam bigblock8.INIT_37 = 256'h34322e06b3897d92d96c4e737c5c677a9c501e5f4a16a372a58e59614f171922;
defparam bigblock8.INIT_38 = 256'h415603abff807274fffb94b9967361842f43dbb714db594acc2ff086fa207b27;
defparam bigblock8.INIT_39 = 256'h4ee362c0210b2418641607ebe073a44f5a67595b304d1969dad2192113ea99e9;
defparam bigblock8.INIT_3A = 256'h03b46e1209a8623c1e5a1ddb2b3c00ede070a4200e63c8c0edb199828ddebe75;
defparam bigblock8.INIT_3B = 256'hffdff9dedfb78e0584478e71d94e5b08de74df347debcbadb77a83309405f34f;
defparam bigblock8.INIT_3C = 256'hffdff9d7be7fd35a5ffcf9ff39cf56ff0ef389768fa7db7135493fd73ebea671;
defparam bigblock8.INIT_3D = 256'hc8e33d3bca319eedd0daa623d3902f123e6e0a61d3a7ffff0aaaae9c89793fbc;
defparam bigblock8.INIT_3E = 256'h915f570e7169a5a3cafb98a539ae8e9e8021c09ac6012c2d5f14095e11e518f6;
defparam bigblock8.INIT_3F = 256'h44dafb057d938f8381c02347f2ae6c5b48500000d51062703695cc12ab83bc5e;
defparam bigblock9.INIT_00 = 256'h97ddeeded68d73f7c562223d481417ad589c281ac401d52acf59597949026bb9;
defparam bigblock9.INIT_01 = 256'h5ca5571ae2127ad1b874d4305db1fbb21565b513648cf29fbd596940e798771e;
defparam bigblock9.INIT_02 = 256'h1ec1800a15613e55040eff807274fffb2e5bd2cbf6024fcf91e786863840036c;
defparam bigblock9.INIT_03 = 256'hc3f446d1470f4f586d5acce4f0008b1e0f2a091587805459898d0056a63cdaa2;
defparam bigblock9.INIT_04 = 256'h9bf32382d3113d9ef6ebee6215b6be69b5faa41f55d755dfc3b1e0ac35a57eb3;
defparam bigblock9.INIT_05 = 256'h5750406604c7190fffae55ff8815d85b1e152d29998d5a99aced8b9076ac32b9;
defparam bigblock9.INIT_06 = 256'h7ab60cd86d099fbe1895128a30ff7d916ab2056466270a1f362a543a302a788c;
defparam bigblock9.INIT_07 = 256'h953d392d0c7aeb0e8935661d03e513af0d407439618f201192c661d1fc57d6ca;
defparam bigblock9.INIT_08 = 256'h2d6dbc5769ffca65158a03156be2a3363d3955c114b48c0eabd7fd0d36235c8c;
defparam bigblock9.INIT_09 = 256'h73ef38d6dedfbd9e8c413d7349f1f17e1158aded3f76d36e6b6f3cb06df68d99;
defparam bigblock9.INIT_0A = 256'hb4ffcd7cde3f1e9ad7ffef5abfff19cfd79799f8bb6677f1fffd6f22ba6b4ff5;
defparam bigblock9.INIT_0B = 256'h9deb1b17239e4a2110523ca9b8ac45241555d5ccd12801ba533b5e35ff1f5f76;
defparam bigblock9.INIT_0C = 256'h0010c4a4cb0235c3800216616358051dbd807074fffb276a4e342d15102a6039;
defparam bigblock9.INIT_0D = 256'h00281840d351252cc994412acbfd803427a690000b928b6c08988780603db157;
defparam bigblock9.INIT_0E = 256'h1b8c656e7f1314dffc8e0b375ba468da2e6c0e67b50829f9aec9432d7bae0396;
defparam bigblock9.INIT_0F = 256'h51b7e623f75e28265fde704ae8cfa1c6c8017c44243132204687e16ebef8113a;
defparam bigblock9.INIT_10 = 256'h0c2c0194347f644f4309949ba7eb47620bff383f12e323d9eedb8d7aeed2e28d;
defparam bigblock9.INIT_11 = 256'h9802544c0222822f45233955998bb33f488ad63c547cfade1086ccf68db4a8e3;
defparam bigblock9.INIT_12 = 256'h69adff845e11ef76ea62bc51a91c4229090113aa688e71b8cb8fcb4b78eb4dde;
defparam bigblock9.INIT_13 = 256'h64fcdd6ce31ffcfa23b3a78a953782eaeb3d0913bd078d9f1d23bf92ca0e4989;
defparam bigblock9.INIT_14 = 256'h426e128c98109d7c5bb5f9c2a8cb7ff50331e7eddd68fe7e939fa92a1ffea7f0;
defparam bigblock9.INIT_15 = 256'ha12386da07d2000b6080470c2ecd6f737f5cad6e7ec483e3b637729d4f6e48db;
defparam bigblock9.INIT_16 = 256'h70c8a61835770c3d251abd0102db8a1e232e5de9204b80037485fb726bff1141;
defparam bigblock9.INIT_17 = 256'h9ee3c25c98f89a7de4d5084100ce7f3be244e1880a3558c468f0030c6ee8648b;
defparam bigblock9.INIT_18 = 256'hd6cac95d1790670792ba228531de7cb2921716a651a60bb674f422b7ae62cc3a;
defparam bigblock9.INIT_19 = 256'h6e471889d5f4f6249171642a9d964eaba6fb767b9c8ba4998fd75d8c45f5df51;
defparam bigblock9.INIT_1A = 256'hd72531a5cb0806b20010a10d380a034f8896fbab7255bb45751be84504121bbe;
defparam bigblock9.INIT_1B = 256'hcf4cf72971378c1b10d0a0449adc289afeb8da7f362ce44ecbab926123845dcd;
defparam bigblock9.INIT_1C = 256'hfccb767f932966bbdab90720185450e39b9041f4a10cb3ee1ab969e9fc1b7395;
defparam bigblock9.INIT_1D = 256'h10c9a5f3723782dc18226ae0479d8b0116145d1692d9ced9a659a0e501193e43;
defparam bigblock9.INIT_1E = 256'h2436f5b4673ce365a1a151e7004fc000db42ce8aa9742a796155214d835ddc7f;
defparam bigblock9.INIT_1F = 256'hfb7223ff59ad31b78e26714408aa666787436448940baae7c96152e0acbfd32f;
defparam bigblock9.INIT_20 = 256'h130caea8668a16e04499e1754c582302a700c23b0a16c82fdd38175b00037492;
defparam bigblock9.INIT_21 = 256'ha1f165a7fbfed5fc2f104fea002ef42be2cc6cee34ecb8e21f99310d4463a13b;
defparam bigblock9.INIT_22 = 256'hb4db9202399dc1f4aae4923780dc323fda8b174e7faad36e11fada69f4274d1b;
defparam bigblock9.INIT_23 = 256'h68e58f4250b068971521cba04d26584a053c0000a608c812040e9d338a0c823a;
defparam bigblock9.INIT_24 = 256'h590f245a544f2ba2ba9bd7cac80f314d01f78e573f1c3c603ee54f19879d1488;
defparam bigblock9.INIT_25 = 256'h9a80825eb19c1c74eb934161a5ffd57f05a8e9c4167b330c0b63f8d297618c77;
defparam bigblock9.INIT_26 = 256'h03e6d503554ce9cd99d1ce05857a650f7dc6b8e30011040093d0b2c0ec94cfd9;
defparam bigblock9.INIT_27 = 256'h31eb6738ea512eeb6946e4af312a2a120d484c915c0c026794405404d8d66f85;
defparam bigblock9.INIT_28 = 256'h5ccaad6d5c11b65b0fe072916f980a476d9d0e963840c02c8ae06d118904330b;
defparam bigblock9.INIT_29 = 256'hf95f000274a2fb72efff7568df0f3e15c8acc36ab7b4d3f5effe33edbec1aab2;
defparam bigblock9.INIT_2A = 256'hea17cff769fe130cade86c8ab6c0e498f96e0ba4030c7301a23bd018862c5bb9;
defparam bigblock9.INIT_2B = 256'h8635d9d028165890c786f45e2ad88f4737d25ef6643408e9371b4161004299ac;
defparam bigblock9.INIT_2C = 256'hce43b4853e41c1ca5192ec0c991243a21869070ee6cac0e54949cc0c68cfb1c0;
defparam bigblock9.INIT_2D = 256'ha4954ffa6f560904cc15a339d9ea0487423a95e9b7c4418a7c86b93671a52a57;
defparam bigblock9.INIT_2E = 256'h91b9a4db000480829c8b2e6124cf4f339eba3f622c142b0fcff4b7d6866a57b1;
defparam bigblock9.INIT_2F = 256'h58cf208c3259c5073bf64f3beeeaaa0e840a76903e845a3af953b6b174213035;
defparam bigblock9.INIT_30 = 256'he4cabc974c08112cc48588f8795b244863909eda8f1acb849b042d1420c88350;
defparam bigblock9.INIT_31 = 256'h5bf97a06a9931fdc6acc955987ddee2c8d6c5cdcfcb44ca64b329908d1eb5f2b;
defparam bigblock9.INIT_32 = 256'h61aadb786dd63651be681d9e0fc145446766206316aee33464feb279d057fbeb;
defparam bigblock9.INIT_33 = 256'h2a22c316ddd0d44d000274b5fb7070ff5a0b454e236538883772a0c59c41e4c2;
defparam bigblock9.INIT_34 = 256'hdd916c1b5a95dd845ca8606830886ef4a594584043140b770a79622cba04629b;
defparam bigblock9.INIT_35 = 256'h028932413c5e66706c1d34592ab7551f0548845212e9994c473c42ec047b12ca;
defparam bigblock9.INIT_36 = 256'hbb469c2cd12961a15be7a2ac4f6cd8627d858c776d65247a8b38b7166225546e;
defparam bigblock9.INIT_37 = 256'h6fb338dbde4d003153babe9fea1812d53665978b32c567a1320db7abf9ea0adb;
defparam bigblock9.INIT_38 = 256'h03eb5535baa9ec5a7995fcf70f3702155d8dda6cc11d9c03f18254645b5b5905;
defparam bigblock9.INIT_39 = 256'hfef148ea2c5a46944df41115798dd922dbea4a511572fa4020389692d4686c12;
defparam bigblock9.INIT_3A = 256'h9b55cfcb2641fc907a9d12675975fbf3e201ed15ca1bfea0cd32c78d09448092;
defparam bigblock9.INIT_3B = 256'hdd1552c12a74202eda9238db9b4e9fbef572f5913635d69655d6dacdfad50b13;
defparam bigblock9.INIT_3C = 256'h69ddb45d024426d8a0671e6176112cafaf128ebbd93e78c6940796a584b69e8a;
defparam bigblock9.INIT_3D = 256'h060a00621bca2a452f0868c9425e02afc2807274fffb04917712806c140f0c4b;
defparam bigblock9.INIT_3E = 256'h71cd41fb83561ea6b4790b58f11aab32dda99d382821136fa09f24ab794364dd;
defparam bigblock9.INIT_3F = 256'h000ca761beb838161d939fc847292c70bad9e55bffdafd4b2d6326f44dff872f;
defparam bigblockA.INIT_00 = 256'h36df2b9a342537e3f866e4ce5a0c796ed866c45eff687d59a9bbd5efdea8c3af;
defparam bigblockA.INIT_01 = 256'h59e749c1a7567f75b3ee03b066a81dda2b32aaa3f747fa945f376381d260c78d;
defparam bigblockA.INIT_02 = 256'hcd2a16de5d6c2a6bb54d91eb16c741629f124f88da0124b4368a124ac286ead5;
defparam bigblockA.INIT_03 = 256'hfcb280ccca51f7ff2c9c36573bb6791be6fe194800e780a3e3dc15e52624ccb7;
defparam bigblockA.INIT_04 = 256'hc89ebabef9f339d4cab41f79f6f483ca7dd485250dfe3f512995adf68809b1d2;
defparam bigblockA.INIT_05 = 256'h500dfaf245b208888d1fcbed18c016d46d55475b522692046fc34324796615fc;
defparam bigblockA.INIT_06 = 256'h0a2e0003469e89232f983688cb4e5194c91a68b1d08a1ddaebd45109966f94ae;
defparam bigblockA.INIT_07 = 256'h18b875a67907088b0105ec2a2884432868c92d5e027cd0007274fffb80a65d77;
defparam bigblockA.INIT_08 = 256'h63a5830c0ecddba315ccb42dfb1bd516c8cb2ecd720577f221f1b461136f80b5;
defparam bigblockA.INIT_09 = 256'h5550d022289e6f767a70fbe5c7fb3b7f6ffafff48dfebd0a03d9c23e889796d2;
defparam bigblockA.INIT_0A = 256'h284757ed214c557e9755523532d833c4f3986bb54723519289a4ce11c1811921;
defparam bigblockA.INIT_0B = 256'he4fe5d852f13e0696138b1d23bfe90002008c6992a42a400013eccf9ef2e5b1f;
defparam bigblockA.INIT_0C = 256'habfb850b0a5ba1712c8a31c3ba4ab86829077fa33b5f64bd6aa2fad7af65fa2a;
defparam bigblockA.INIT_0D = 256'hc51671d7aa872080a0d6ec8bfa3e23e9ffb3d3d1e31fa9bfedfa18347a7bddc3;
defparam bigblockA.INIT_0E = 256'h51d99ccb2255ae86a559214f08db94a10ccd4f88887746d7226eb6881f87c959;
defparam bigblockA.INIT_0F = 256'h4336241d8442213cc8101c554890e30265a8e1f880ec06feaca696c030992c4f;
defparam bigblockA.INIT_10 = 256'hfffb47570827d3c2e3c12b8822da71d7399bf9706d9b272583ecb0b61031186d;
defparam bigblockA.INIT_11 = 256'hb41390ef209824567da335330c4a0062dbed280415ba6926585e0312da807274;
defparam bigblockA.INIT_12 = 256'h0495e6aa4e8e7d3f7f64ed3307efbf7dfeb11811aa8d4eed8be04b78c2600858;
defparam bigblockA.INIT_13 = 256'h5bf40d3454428374b683eedf0bb80b12686edafc2ec60248d400f5002d9dd03f;
defparam bigblockA.INIT_14 = 256'hc5388980a1a0e50f488117040220cb3319e5dd4cdc901adfdb0aa5a2f5f9dea5;
defparam bigblockA.INIT_15 = 256'h341232feb9a5d4f1559998e368e72d9e2bb1fdb47b63fc4fe0843c90824d8951;
defparam bigblockA.INIT_16 = 256'h46bf29b70c315f33879e475f1aee23ead58dfa02a434cc0296ad47e6d630efe3;
defparam bigblockA.INIT_17 = 256'ha03db100291791d5bb2d566ae39f0a0d89e5b565118d8022cf5c3f663a755b46;
defparam bigblockA.INIT_18 = 256'h178dc29640e2a0468848407320955d81dd8116fbf121d43af52c10f4884a4f72;
defparam bigblockA.INIT_19 = 256'ha9e31876ec4956b3e7dcd42dc04753b89d5bcf4c999a80b75427dcc7a1388cd8;
defparam bigblockA.INIT_1A = 256'h02c1e4807074fffb0da59e169a313d5d8c183db7301c41de74f9f1f0b789e225;
defparam bigblockA.INIT_1B = 256'h89fa1fa119b8b481946ee0af945875445535080a01221baa2b652bc8698b4d5d;
defparam bigblockA.INIT_1C = 256'hb69f2512ea1a99951ea1f56be10bffff12ec00009ff5e06f22ca5ddb48223052;
defparam bigblockA.INIT_1D = 256'h05e6dde3000644801282683fefcbe221b6e5f5104d466aedbb44f6edf614b436;
defparam bigblockA.INIT_1E = 256'h93f6850091e9d68b491fb5469efa467253a766e37aa3a584e8a1431ba477d150;
defparam bigblockA.INIT_1F = 256'h2fd9ac47a4e6ae794169fe712a236b38e6ed5d83ba90086f7dbd9bb975ea98fd;
defparam bigblockA.INIT_20 = 256'he917ffa20817ff20ffffffffffffbffffe9a05907774e5f7dcb665dada3f3d3f;
defparam bigblockA.INIT_21 = 256'hd401186a8554dd1db7b8ff2f465e263dc8f3af4124d85a619c511a4ea31b0348;
defparam bigblockA.INIT_22 = 256'haa5d36659e127ab05dc6e2eb46796c36c8ddce0796706f0bb13111cfab1344cb;
defparam bigblockA.INIT_23 = 256'hf0e27f58848795045e622f43906030d2cad7728609bad48aefc9c62c1764dae2;
defparam bigblockA.INIT_24 = 256'h3829272e5bb1b64d000274eefb72fbff6f722c6ffcf61f55554f674909d3ba23;
defparam bigblockA.INIT_25 = 256'h8d77009b004053e88e7e38b293156de4ab94ba60c49c096e4ad1050e7701e4db;
defparam bigblockA.INIT_26 = 256'h71d02f2330fd53a7d3e7f91f657a7432219b5961ef0747be4fb90c76f0f472f2;
defparam bigblockA.INIT_27 = 256'h2bd5d818eb6506809cb4579670c2a69c11fd588e346c2d1f019c19500200c3b2;
defparam bigblockA.INIT_28 = 256'hdf7677c7ac28a57364ceaba2d41feb530e73f4e10eff44c63768773e581e7ebd;
defparam bigblockA.INIT_29 = 256'h5ffebe8f39da7548c1b12d6b30b753f6dc216d9e7602170990d2ec5026d42c1b;
defparam bigblockA.INIT_2A = 256'h6e47282d7711d9d0f9038b18a8cded0bfcf6fff04a8938b12ea51ae401490801;
defparam bigblockA.INIT_2B = 256'h70a381f3384f45492a4ecb9783630a4802ca400172a04c876f17e5e7b7b6dcb5;
defparam bigblockA.INIT_2C = 256'h9e6b689b45722d1a90beeebcfc8689a61b7cb9acf7d46152b9dd942b369b8a90;
defparam bigblockA.INIT_2D = 256'h29bfa9e528ff971f9c6d109b9994e39c5b62a4f1c83f2009f368bf42890b3587;
defparam bigblockA.INIT_2E = 256'hc20e660044dbb8258b54db391047000374f8fb72ccff6cafd27ba617ac3ea8c5;
defparam bigblockA.INIT_2F = 256'h8d6748d2034c19d1c63d36d70a0a04001980619e6d9ca013fa60a6141f6c0af9;
defparam bigblockA.INIT_30 = 256'h00130402062933947fb8bd4d9e7e9dfab323da837261289e47ba9e1e7e210a67;
defparam bigblockA.INIT_31 = 256'h96231af9f5223f9798cae24861a8a213359ef6c570ac7c7e17ba519581ad75c5;
defparam bigblockA.INIT_32 = 256'h5453f59874e64060b3cd3f514171b69d792dcd5efa3513a027163199fc274358;
defparam bigblockA.INIT_33 = 256'h28e34020ffc0d5ff6ebb3147876717959fe89a0218bf6ac28365007661769c41;
defparam bigblockA.INIT_34 = 256'h8e90feaf3bd9009f00bc64c528dbb48b35554f8b9a1d8c2b01c84a2710d35db6;
defparam bigblockA.INIT_35 = 256'h243d790f624ae4c73ae43aa363e364a319aac905a4ae0400a801c1dc9dc4995c;
defparam bigblockA.INIT_36 = 256'he27f219a8d64809eeebc0593b38a00c6bc08906d28c6e7ebf58a8647aadd6d2a;
defparam bigblockA.INIT_37 = 256'h1c4fad669bc98c7dfa0fa59b59fac48bea881e50b1fa709cfe446e2f50603197;
defparam bigblockA.INIT_38 = 256'hc4a01d6a0bf9270e5701851ba82b8716dac9ef46800274fffb7200ff53fd15d1;
defparam bigblockA.INIT_39 = 256'ha5d121c572b9ef79d54f992fe8dc890431825dd3a36d609262a26d68b393f8a0;
defparam bigblockA.INIT_3A = 256'h0bc9279cb45a0cb00490103050af292837aef8612ee8dbb3b584a703aca2c326;
defparam bigblockA.INIT_3B = 256'h70e7053fb7bd35beeed15c12869d4c6e6a5fe168ad7cb41465fb6de56a09e281;
defparam bigblockA.INIT_3C = 256'hbfa477fd9cc31f2669ffe503ce2d83e7938a6ad27ca5657c8d33f8e00d1ce837;
defparam bigblockA.INIT_3D = 256'h216a559e830b248ed669425c5b47577e71b82004e020ffffffffecf4efaf1bbc;
defparam bigblockA.INIT_3E = 256'h4a6405222001dbd2df408cd747cac7a7f1fd0c4d8e267920b67fd72a6fb8a292;
defparam bigblockA.INIT_3F = 256'h00b59be67426162293d6c26f5d4549b4c2f8a2a5bc366c5cda15bcfc85d7e594;
defparam bigblockB.INIT_00 = 256'h48c8cf6326bac5625d513752da1c9ea7226d3e40e7a92191c4d6391d5be48009;
defparam bigblockB.INIT_01 = 256'h00ff800825bec8abcb12444df7cd7457c24bde71a9975931663a301427361a5d;
defparam bigblockB.INIT_02 = 256'h6d4cb2945660c6191d6a0bb967785718651b382b8a16dab1fa47800274fffb70;
defparam bigblockB.INIT_03 = 256'h50193753e14b36956759050710cf1404921d02af5c6559741af700b728099116;
defparam bigblockB.INIT_04 = 256'h7314cff593eeb2328a702486a167a78d95578a10622a124ac9d0b3b64b74904b;
defparam bigblockB.INIT_05 = 256'h048eed82d4e582a8d027dc7c13a8ef9774175a8522e1ec79cee13f2c9b381330;
defparam bigblockB.INIT_06 = 256'h7fa6852bfce2cbfce7df6a32c2fb4c6da5af9d0a1bddf881a35700f4ddeb0c79;
defparam bigblockB.INIT_07 = 256'hff86e2efdd378e93f8f49b5e6b3affebe3760c6bda625f5bcdab297bfc5d358c;
defparam bigblockB.INIT_08 = 256'h50d8b19e2606252c5c6a18b26443ed1dae4046dac00099f4a6bffd76e7efa8ff;
defparam bigblockB.INIT_09 = 256'hd5bccffa93fd7ce9656d4d09c4a08ad79bdfeec1a97b2b901f919b6a04ce0cef;
defparam bigblockB.INIT_0A = 256'h04a91157e49758bbf578d0b130b968c4d4ad75279c8c4e8891e500000000535f;
defparam bigblockB.INIT_0B = 256'h02abff807274fffb2b0a95d32b221711c689759eb1588ea3c54e8290da5a10f1;
defparam bigblockB.INIT_0C = 256'h8b4b1cb615682894136d20ba255168465537c00c2447db472f841630318741da;
defparam bigblockB.INIT_0D = 256'h2e5c84315d92d572d0f79521d8356f8f144d30dc0d51cefe895fa6a67c6591c7;
defparam bigblockB.INIT_0E = 256'hfdadf4791af77de76d668ac1816c2469110eb8231dcfeedb67c7edd355b810c2;
defparam bigblockB.INIT_0F = 256'h1fffe0e00b83e800fd16bae583ae18ba07f0fffeffbf7f07727fb0647162cb82;
defparam bigblockB.INIT_10 = 256'h5299d133c735948d1c1851fa2ac525d74cace54085225dd0c2ded12ec24bffff;
defparam bigblockB.INIT_11 = 256'h59ca5bb8a8745b2db496ca6e91560913f33de4e0e96c22d1f12432c397c769b3;
defparam bigblockB.INIT_12 = 256'h1f0e19ad1ca82c3ec25c0e9bf8623ec1d990783db72d95c0a854bcfa84ec7242;
defparam bigblockB.INIT_13 = 256'h1edcea963d5e253a2e5e67b2172f72ac36d19e9cf2cadea19350075279069f40;
defparam bigblockB.INIT_14 = 256'hb5acf6e5448e8eb54abe2a27b454e78cc95fc7482a14b321ada276b0403bf04e;
defparam bigblockB.INIT_15 = 256'he008853d4cd803daff807274fffb3fecba6fbd2b516e71fab547f50d72965aed;
defparam bigblockB.INIT_16 = 256'h7bf9d7ac9bb95e66396ac0004b1e8f2c00f587806259ed190052a624db133804;
defparam bigblockB.INIT_17 = 256'hffff0080ff00dfcea266497f666b7d2663ebf46a66fdffa68d6da6d2ff36065a;
defparam bigblockB.INIT_18 = 256'hd68d1a9c6e6c7695d87d445648d17998309117402f2dd324330662237260fffe;
defparam bigblockB.INIT_19 = 256'h9fd565bdab446915a714cf544bc0000d204014d0129c228e455f55d7f5b44156;
defparam bigblockB.INIT_1A = 256'h9dab0b60cb554b31189c800b5912bd9d92aef7c689c7ed909eb03221cf509603;
defparam bigblockB.INIT_1B = 256'h1da19d2c0fd261741b0146fcc4b5d99a45e0e2574757af374ba8b197bd47fadb;
defparam bigblockB.INIT_1C = 256'h1e8ee77a5fe874bd3fa7b177e6f73aa4ee528fec8da3639012204fd66df7149a;
defparam bigblockB.INIT_1D = 256'h1fffc0804c636633b3b1e4de5dbaa6e6d4ed7a69fe98dd7cede6696bf48ef93d;
defparam bigblockB.INIT_1E = 256'ha582109d56fdb1e67ef805ab7e6afd3fbd5b909459a221d843a15255d933cf07;
defparam bigblockB.INIT_1F = 256'hc624cb46328380000661645a04e0c6807274fffb0864ec42e41e2935b8485475;
defparam bigblockB.INIT_20 = 256'h6447ef55f72459619419cd6446b0e86e90011b900b6d208bf60068dcd9830011;
defparam bigblockB.INIT_21 = 256'h1cbd47b97db5a32e91f5a9003779144b2a9c69b1b4bba0f7f4e0355c8e612372;
defparam bigblockB.INIT_22 = 256'h40bcdeba57ab2b27ddfff79d3bd9066e15d069cea73f80145b25573bdafe8fa8;
defparam bigblockB.INIT_23 = 256'h991a22446016d50cdc6bb33ab6170c4c7f0975345faadb44d8e1f74cb4d6e46d;
defparam bigblockB.INIT_24 = 256'hbf1c981c07a39fd3f9900c8f368a0c1f30b9156c3a46a55348126a4245406536;
defparam bigblockB.INIT_25 = 256'hcaeb59aaae6556a951ee59244a54ea9e9a03de314adf9a20959a0248503d8b3d;
defparam bigblockB.INIT_26 = 256'h0439e8610969d1102a26a2a24a48342736360a0b439b3abc6865bbe5f79432cb;
defparam bigblockB.INIT_27 = 256'h2652ab706fad9e0ce0518e8fccf373d059cf1e09b3871480c7dd209b255f236d;
defparam bigblockB.INIT_28 = 256'hb87f521dddcb722586afd32f044d562468fb09bbab95a28860ca4ad5532e2d4f;
defparam bigblockB.INIT_29 = 256'h75a34d072c4c04651ba71b831622512341dd02dc91807074fffbebdaca2d5b0e;
defparam bigblockB.INIT_2A = 256'he6e6a596efbf727a48ad6581d0c8821d9b5eb2799fec99d0a8518dee40822055;
defparam bigblockB.INIT_2B = 256'h28640e1557657e930c28d5bf5dfc91374a9f0be3fda33212f5b34368faea3a99;
defparam bigblockB.INIT_2C = 256'hbfb5acbed40fd7125bd7925e902342db8b705cef63b704e94909c8db062f6288;
defparam bigblockB.INIT_2D = 256'h46d793f345868719cc28090fd8bda98e3da74e28889ceba7a180451236b42c50;
defparam bigblockB.INIT_2E = 256'h49874f9308c8bbf7abf0480eeafff556f7ab6e6afe8502591dc9a80f00859239;
defparam bigblockB.INIT_2F = 256'h734a0d87d53bc546d3c2a235449fa262b93ae95c6843ffb924f552e776de56d6;
defparam bigblockB.INIT_30 = 256'h10c42beb2cfa299caabc70078f9cb3621afd9148161617832b9a1b6d7b5934c2;
defparam bigblockB.INIT_31 = 256'ha0f89acfa475644c3a0b33f0bc956939c156a8cd8c6aa15218a8002024820401;
defparam bigblockB.INIT_32 = 256'hb9ff31ee761e9f4068b9846de4cf4f3fb71195e6ea28f2b7e1560550d58cae1e;
defparam bigblockB.INIT_33 = 256'hefb4830d6fe0a6200b790bf12874ef18e2db2220cc2dde68e7470002749ffb72;
defparam bigblockB.INIT_34 = 256'h53debca4d727f2bc4a69452b94569a1c25be6fde6bcdcbd7710a97d808823095;
defparam bigblockB.INIT_35 = 256'hee316f0c72b4509194363af7554c8ce56d04c923000d018049e12d09d0e24769;
defparam bigblockB.INIT_36 = 256'h71b713d67b0a3e9edd19b0ef585c4c1a59611e10c1b7890b42921b2001994400;
defparam bigblockB.INIT_37 = 256'he3ea0fea1351256aa41404fae691ae58a3e777d17e9c92aa93ebbe50ce23605e;
defparam bigblockB.INIT_38 = 256'h0200086bb1615448709cb51eafd463a141e1c6847eb2d0e3236f4dfe9a366444;
defparam bigblockB.INIT_39 = 256'h100004006b08f983af044fbc0b1a955f71a70ad79f5189953583a7638db414d3;
defparam bigblockB.INIT_3A = 256'h9bff5dfbc6423f9d294a4c45a3845939422a3686d0385dc8688c8e502da425d8;
defparam bigblockB.INIT_3B = 256'hb57f74ca22f57f90345d1b7ed87fbf54006ab180be835c7241dd2b11a8482447;
defparam bigblockB.INIT_3C = 256'h000374abfb7200ff56420045ebc467b4d16965249d079b55dd15e9faf5abfabf;
defparam bigblockB.INIT_3D = 256'h05724800238a6e28750cb6e044a00b710c1d63068d0ca1cb2a15272edc69225d;
defparam bigblockB.INIT_3E = 256'h3735cfac8c6efda7b5601d850000491981c607becb9435648424c830495136dc;
defparam bigblockB.INIT_3F = 256'h716ace83608c2ca28608568aed68475b904be39014671fce02ce44b3e0e4bc2b;
defparam bigblockC.INIT_00 = 256'h70e9479fc5da5c54b5b6f9e2d1cd94407cae6660cc0fd4b2c9b680802389bcf4;
defparam bigblockC.INIT_01 = 256'h00008800ee1ec1e792edffa2ef3fe62f0879c3651ec559ce6bed7ddaffc5ff93;
defparam bigblockC.INIT_02 = 256'h96a352243d64436549b620899188e5a9bed1f9a351aa32060c83459c2369b249;
defparam bigblockC.INIT_03 = 256'hbe154e3a7e759a4cd82ffab7c1b7f56370d7932e41c962c339f14598ae3e5dd7;
defparam bigblockC.INIT_04 = 256'h54bad49fe7ff28fb6459918562dda86c63d8507e0eb34bd0d9d517ab3f84a8fe;
defparam bigblockC.INIT_05 = 256'hc88146daa59220a0b10802104c94a40928b95fcc4acb49707b76cab4bd2821e4;
defparam bigblockC.INIT_06 = 256'h2c2b5ad1df4f000274bafb72c1ff600deeb73105a7f8d7a0628e39306d9b2a54;
defparam bigblockC.INIT_07 = 256'h49cca6105229a4a0904a63986d745b0678e8c61d0d6a4d6d23505d20017b5016;
defparam bigblockC.INIT_08 = 256'h286bd49ecb943efc9538c79362589136995cb58b5d02bc0f7aaa4716c1ba84ed;
defparam bigblockC.INIT_09 = 256'h9b65fd29badfe4b4244d4ca065f850cd9ecfc2d9b39406f7350a7ad1c68f1037;
defparam bigblockC.INIT_0A = 256'h3e716da546a39c1d1ec7cfda98e4a101cd55994008c23997ba50353dc9bff0f4;
defparam bigblockC.INIT_0B = 256'h911233881b284e644249e4012285c2f0c86404876f624a04c65b989fa0c94327;
defparam bigblockC.INIT_0C = 256'hb1b1a1e37a5ee837a3c469001327a46e67e8b4c5631406ef2ff2414c2160931e;
defparam bigblockC.INIT_0D = 256'h990ad80c290ea72753f45cae182f7e628dad14f5aae23ca267bfa00e302ec752;
defparam bigblockC.INIT_0E = 256'hdb558d24808a0188daf2549a02d640be06f695d66ebeefd80830fabf658e9727;
defparam bigblockC.INIT_0F = 256'h85902539800125801a1b4936c33381373eb5d082d0ebfc36286d484691485b1c;
defparam bigblockC.INIT_10 = 256'had0ce2db281d2b3edd69194d000374cbfb708bffd471a996902a688eafac12b6;
defparam bigblockC.INIT_11 = 256'h003b363467466b2ecb8b0de44cb1c0ce308c6ea8700b78a0a49433750be1463c;
defparam bigblockC.INIT_12 = 256'h59f9e5d4eb13be82e5cc7ad685b9a3a985fbb265b7dc16ff9c7302298547062d;
defparam bigblockC.INIT_13 = 256'hf0080ce0f4b854cf7efdcf0ec2b21d929f0193f0cf4ea7be710bfa58214bd91d;
defparam bigblockC.INIT_14 = 256'hfdf6bcd0a8442e740b20002600208124fae169099a97f68776a4df36a77f4400;
defparam bigblockC.INIT_15 = 256'h95ef160466cababdcbb2b70a87739fb467af23abe84be2cc90d6799b745a9132;
defparam bigblockC.INIT_16 = 256'h9a9a0cad65ec23c572fd8b66d59134128430a9bb2899b47666d6cb8a83a72d13;
defparam bigblockC.INIT_17 = 256'h001086ab1872f901d0b0dad32ce803940303c80366428a083c502822562399a0;
defparam bigblockC.INIT_18 = 256'h3606a21123c581aa00010000a98134ff72953b8066d2b686ea2dd5057fff0002;
defparam bigblockC.INIT_19 = 256'hd30cd0863480e0e7cbd4026bc43ae45eda18699255ad11cec96e2b54c7a19caa;
defparam bigblockC.INIT_1A = 256'h71475933580c2066db8d20421eba51224ddc0324d7807274fffba68db391270e;
defparam bigblockC.INIT_1B = 256'h6423233bff241985d98308b7769cac88c9e75101dc418d49306005eee84ea467;
defparam bigblockC.INIT_1C = 256'h2c00c899c423581fda6ddeffd3f94fcfffe7def9579dad8ef72ce9a799a1999a;
defparam bigblockC.INIT_1D = 256'h30764ea02c06012a0000081a828f8992782c167b7a12987d695cb49304510000;
defparam bigblockC.INIT_1E = 256'hb0830c38a6b12114a89038b4e4080d52c2cbe60e48ba1c2cfafa4b8381737ec1;
defparam bigblockC.INIT_1F = 256'h40afc51669c766a49fd2943934e7050ebe9d07f55b8f58a05105dc85355b51dc;
defparam bigblockC.INIT_20 = 256'h4000a0f5daab1fcaef16f133427549abc50485bee9197bf3169166c2a666bc3f;
defparam bigblockC.INIT_21 = 256'hc9eaa866a14cab41000ab800514b67d91b25bc42c358a46814c9dc4a97ff0000;
defparam bigblockC.INIT_22 = 256'hbe84a32957259347d182ae2037597dd53ae1bd531c5a11954244046e41a3c372;
defparam bigblockC.INIT_23 = 256'hcf62a39c383b9fe06ddc46b7c273a7285968b9b4fd7aa8b24e75bd43cfb8c9db;
defparam bigblockC.INIT_24 = 256'h852d285818736ae6f565140c0526ab5c15411e18b18643da0360e5007274fffb;
defparam bigblockC.INIT_25 = 256'h5fca4c26ee7ea7f2588238544c8bd3e229bf3b2c327638b520bc25d220517413;
defparam bigblockC.INIT_26 = 256'h3d706172da4b2a6c707213b628a3b68f1c910037cc00a3f233b6c6174dffd4b8;
defparam bigblockC.INIT_27 = 256'hc800d6e54b49862eaecaac0ee35228543c4c0830b9096d8f05d4920000181b02;
defparam bigblockC.INIT_28 = 256'hdab5b6f6004735812bfbdb4a674c78b6cc7c31e609665a7b70087d41b651dae8;
defparam bigblockC.INIT_29 = 256'h1dc9b132f9f2417e72708cf2615959fe84a47ff961ebf48a2bcf43bdc53f04eb;
defparam bigblockC.INIT_2A = 256'h2a93a287487a19a8143667e8a069e46d049434e00fc3056ca5016513080ac251;
defparam bigblockC.INIT_2B = 256'h1e1bbc253e504d12a924428c1730003a0102a2a05262f39090c67450167d6e41;
defparam bigblockC.INIT_2C = 256'h387cde81f8a76d2185bf6b6c1be68c6073e7f610fb4bd633e6d149d9bb7f9cc0;
defparam bigblockC.INIT_2D = 256'hf0807274fffb4c2116fd88e3fd9c1611dd4e97a599949988cf632f0dea78759a;
defparam bigblockC.INIT_2E = 256'h69f69819681405ad2859147e6a664513000e0426ab5c16611d2ab9864d5a034a;
defparam bigblockC.INIT_2F = 256'h40b407754dbe31ca74aad9b3db4525c81000d4205faf303fabeb4b047522b59c;
defparam bigblockC.INIT_30 = 256'h4a814b64352cd2b268f14361a85d62550101c00041abb50b08656a808febb368;
defparam bigblockC.INIT_31 = 256'h86fdf3924ea35dd1552ebbde9cf13e9bfe70ff89f6d86b6d5933a6bcda8822d2;
defparam bigblockC.INIT_32 = 256'hc750833da2509fbaf7136ae5dc1cbb36510e188269c65aaccc0e540c99cb84b5;
defparam bigblockC.INIT_33 = 256'hc100fffffffffffffd5f4f6fa8351bf7cc8c51a9aee16abe1214ebe73ac9da34;
defparam bigblockC.INIT_34 = 256'hc15205eda060217d9698d9644187806b194e502cc0d300c8e5bdd685db7b2648;
defparam bigblockC.INIT_35 = 256'h98bf7631c4a6e67a8cbcc30a49b5d459024a222bc13ea179338000450028df70;
defparam bigblockC.INIT_36 = 256'h89413dca31f6054c2ce7be33d420397bb432aa2d1a6014e68f67238d421e5b7d;
defparam bigblockC.INIT_37 = 256'h51264ddc0363f7807074fffb96d7e3c6e95bb77952268485d9959dadd0dba774;
defparam bigblockC.INIT_38 = 256'hfa1bad24d42cd647083028138d6e607c99517124910d164b04c5bb871f021f18;
defparam bigblockC.INIT_39 = 256'hcdae04c5d73e3ec99d90709af2ad7c93cf5463328747ab1888e56eadc923e800;
defparam bigblockC.INIT_3A = 256'h79e5d1bc57c748c3568db814c7247cd96864ba509a6b6db11881100406c11f47;
defparam bigblockC.INIT_3B = 256'h26864735d8b7d9d1977f4a4bcde296be3fa46e0bef1e5936e14a12561deccff2;
defparam bigblockC.INIT_3C = 256'h4a0ebee23eac7dfcce19df1bab3fe6f6c6dbebb17b6d734d68efc973c87da19e;
defparam bigblockC.INIT_3D = 256'h9a67625965c7a4d4dbac724800c1fffefffffffffffffffffffff57fd1e974a7;
defparam bigblockC.INIT_3E = 256'hc0b23282549a003682080f40966910e14a3f1371b3c193024f4d821579fef607;
defparam bigblockC.INIT_3F = 256'h37517214cda83616adb5c6d763ae4d5b6addaeaf48f61c7ea7850df4fcfa03f1;
defparam bigblockD.INIT_00 = 256'h0a8e3b50df9ba21fae0cbdcd083556c1e26d091fd58ad7d9ce4a7a442c5b3adf;
defparam bigblockD.INIT_01 = 256'h5730231b4823eb16dac1924d800374fefb72e4ffd38c2e9c38a08fa76d103488;
defparam bigblockD.INIT_02 = 256'h6dcaa92410a0dbe9cfa3aff8ea3e5163b1966d4c8c0df140e6240f6a4b75a346;
defparam bigblockD.INIT_03 = 256'h04400ac8c8e844ba94b12a57e569672993c85a1bd9c3cb343697322a78a86824;
defparam bigblockD.INIT_04 = 256'hb8dce677e4245cbce9938519949512e5813f7703136200e284d9788406209000;
defparam bigblockD.INIT_05 = 256'hb22b201bdbf0c4dd95178a237fa9f7aad9c395d4ddeb52e5d490df9b89136b82;
defparam bigblockD.INIT_06 = 256'h03f6d44e44c9a69e4536c60f5ae371599b8e4b6a5e6f8a21e816c9b1fdcfc61e;
defparam bigblockD.INIT_07 = 256'hf69b58f6ae11f79c5b3d8f1f18080f9961486e6429240008f810bb554ebdfe82;
defparam bigblockD.INIT_08 = 256'hc19d8ea772173584919a0fd6898f0000002c00e00354b39985c2970c53906429;
defparam bigblockD.INIT_09 = 256'hd3b955239713075047711dbd01a25798fe8a1eb454498b4bab04c12f0496b1d4;
defparam bigblockD.INIT_0A = 256'h8c353d2e14a1728a506ddacff35e7bfe0a35e62eb856ac1baf806d4e3fc3fc48;
defparam bigblockD.INIT_0B = 256'h376c4c0d46946724c35bf8238959db416f43800374fffb729affd291409ae74e;
defparam bigblockD.INIT_0C = 256'hcecc238dc8258300df4b478b7a6de4142a1cdce0388e04946d9c900db720c62c;
defparam bigblockD.INIT_0D = 256'h00201ff3cf7db375282e37f90991133d592a139229062ed0091921e060127485;
defparam bigblockD.INIT_0E = 256'h9977efd64869aebddd85e3c7e0512b901937a243951129294ed368ce06eba000;
defparam bigblockD.INIT_0F = 256'h1396f3240d5ce5d7c292a5bdcbce9b1bd678b3ab273ecae54fe395676aa66729;
defparam bigblockD.INIT_10 = 256'hbcbb86faea86032c04de4c95d1185cb4f55ae2f3451fa0639f5bf6fbb4b1d973;
defparam bigblockD.INIT_11 = 256'h7a05e8098e597b9a82341baef6cb383c4d6cfc9691c900a4fc104c1bc30590f8;
defparam bigblockD.INIT_12 = 256'h76e4d10412d3b7269dc0211789d1bc38d4aa257400060010aab21ce2ba637349;
defparam bigblockD.INIT_13 = 256'h5deec192f35dbd53322f8de57f7994cc7e96d0dd7a02bd80d61e6eb5ddf268e6;
defparam bigblockD.INIT_14 = 256'hcda31d2a7a3204496de450e76e483955bb14b13c793528db86e67b2da38862a1;
defparam bigblockD.INIT_15 = 256'h928db1e046240d6d0d31c2766a24433bb8252b45db394543800374fffb72daff;
defparam bigblockD.INIT_16 = 256'hc2eee0bb296692571923900031c867929ae7146cdcdb4835e99f4985609a6d9c;
defparam bigblockD.INIT_17 = 256'h7294903200c4120053a834550b486626c4686ee7aa60c0b1388b23913f9157e8;
defparam bigblockD.INIT_18 = 256'hee13708170feef2bfbfe987fe3bfad1816403f7b283098559218662c2534f3f2;
defparam bigblockD.INIT_19 = 256'ha3bb1060840a2eec40681c03e8281a7bfbf0944ddc1ce25d9f2375b9f3112499;
defparam bigblockD.INIT_1A = 256'h6bde764fced910650408cef54dbb73c25d883bdcc5fcd53ebbbb521fbba7c705;
defparam bigblockD.INIT_1B = 256'hdb4472463aa401447df632721bc1db994509d93a143040188324213ef6bcbb2e;
defparam bigblockD.INIT_1C = 256'hdddeab31febb4961fad5280d005d486488d4c11251102b43fe4d293e2c72a27d;
defparam bigblockD.INIT_1D = 256'hb93e3bbcfee99f05987794f90b41e753716ebfde26c69d5d79ddbdbd2b85530b;
defparam bigblockD.INIT_1E = 256'h74fcfb7045ff3e4ee5b799956f0fbfd8cbb2f33b39319333ccfff48b98eeaf8f;
defparam bigblockD.INIT_1F = 256'hd043c1892d9c840d4de0e625236c0d2122946724435bc8208b2d5b3946438003;
defparam bigblockD.INIT_20 = 256'hbbf2268a3c5c1971b45a5dbceb9c8e8459d7303d62495e3ef7c3e5d2d64eccde;
defparam bigblockD.INIT_21 = 256'h3130012519ba07d46076ae3718d240f91801428bd76b6db6c723aba51c169552;
defparam bigblockD.INIT_22 = 256'h8eac0e35091a5dbb2a81760ddbb930aa51cc8638c71df7e2b5c9f78452e2dbe2;
defparam bigblockD.INIT_23 = 256'hf7ff9145b4213b14fb5e67b13159da2457d1e287b3be37207d983c918902e81d;
defparam bigblockD.INIT_24 = 256'h01622d5fa29876df4a3f37fddc75936e415711ead317ec650d61dabf76cffd54;
defparam bigblockD.INIT_25 = 256'h45047190cef4258029f326463f1f2b826ab3f22da48a25e1da356da527230001;
defparam bigblockD.INIT_26 = 256'h0477119cdda2dd20e73063a18378c6b1f3d7ad591cc0274baf8a40008235360e;
defparam bigblockD.INIT_27 = 256'hac8ae6b625e15b1a03fe4a593ea0f16dc58fad26695f9c374e614144b1809032;
defparam bigblockD.INIT_28 = 256'hd18860de0414fd807274fffbe84fc316f415352f1fcf3175239536319d1ffe73;
defparam bigblockD.INIT_29 = 256'h87dc2ec28235a9b90c58741306afe055b0c17ba75583020e04264bdd14a14e5c;
defparam bigblockD.INIT_2A = 256'heb8a9bada32b556a0352bc71f4f635ff1000acb8bb2615026fdee543d4c37db2;
defparam bigblockD.INIT_2B = 256'h72d547e9cddb10f3bc2ab1712c32ad51c23a0022dd381fa9d0a8105443eea292;
defparam bigblockD.INIT_2C = 256'h3048e1c039d7d21cefc57f8511070a0bc88503ac81bbae7b99b34db6c77c52de;
defparam bigblockD.INIT_2D = 256'h2623f94335637969f94ae53849b9d8b4b882f9f35c77c68e664b00c46a84534c;
defparam bigblockD.INIT_2E = 256'h99dc8db602a4af8819327d88d72db9fc5f33b65fb6490ee6e26cf31511b9ce11;
defparam bigblockD.INIT_2F = 256'h000010027002f574ac1b69daf2187823189959c82fee747aca04587940baf4e6;
defparam bigblockD.INIT_30 = 256'h7ceb6cedd91213022a83d46585b642ea845508267c870616640fc81a30f30311;
defparam bigblockD.INIT_31 = 256'h1a9aeec3ebec04ba1fd71ff78113eb8d367111b995ebf18f8f5512a1377b8d18;
defparam bigblockD.INIT_32 = 256'h5b9d22e31dc2d1854cdc0330f9007274fffbd8c5c4377b5b1d2ddecee56ee9d5;
defparam bigblockD.INIT_33 = 256'h58562358074ba7fdf17f870137a1141964038c6e6875207573261939160d0582;
defparam bigblockD.INIT_34 = 256'h93bcdb578383edbd8eaa91b438dc3800321cb3dfc999cc672ea6cfbd6b3caf33;
defparam bigblockD.INIT_35 = 256'hb8a403ad120c3d5a5741485012263408226822136e01009d04000300cdc61fe3;
defparam bigblockD.INIT_36 = 256'h9bdb5cbb14d3f989709bd9b17aa26465998259414b296d56b62d67be757bb5b9;
defparam bigblockD.INIT_37 = 256'h860edc95541299b9dca94e878d45b530d35f8bdc93a300332db0dbbe46b40056;
defparam bigblockD.INIT_38 = 256'hec2e73b11a4d72496000d8b08cc5412fc6579b6afb3e7a35c913854a919cde5a;
defparam bigblockD.INIT_39 = 256'ha887224641e19585001414093090d41c445540ac19f29e85f47f965dd33d0d39;
defparam bigblockD.INIT_3A = 256'hfcc13bb45b318bfe95a365876425ad7d48dd96496da1d480dd219223c2d22181;
defparam bigblockD.INIT_3B = 256'h9174f371d194dd1027c8bab822dbd58e5fbca82884377751b382405d5b34587e;
defparam bigblockD.INIT_3C = 256'h29835c0e18665b7721631e4a91885edb0371fc807274fffb52927cc3be96a501;
defparam bigblockD.INIT_3D = 256'ha8522491000716e52d902ee2bb9e7dfcea5be58f8830e814066d2051ac796f84;
defparam bigblockD.INIT_3E = 256'h366406ac00023000c34791606cda4a36f127f68e724932b30f53c889e607674c;
defparam bigblockD.INIT_3F = 256'ha1e133f85b0b52071d47ce3d525c845c3951b421d608314982a138491440f473;
defparam bigblockE.INIT_00 = 256'ha841e5057a735f62596db0a4e4d4887a30cf6a0cf9c100c96e71d8c2c0c94f3c;
defparam bigblockE.INIT_01 = 256'hffe2ffffffffffffffffffff9fff4136f6d1b7a8eb675beff6e87f576c67b6bc;
defparam bigblockE.INIT_02 = 256'h840006d1547f064f995504e7965f8c43562df2cb0484c542531daa4d24711007;
defparam bigblockE.INIT_03 = 256'h0b4384a9988ab1a460c1a20fa43014d429a413a1ba331a95101f9a4ea1380921;
defparam bigblockE.INIT_04 = 256'hb6137f8f0e92df3e655a71217b86076f5f8d90359314430125f42a268f544aa0;
defparam bigblockE.INIT_05 = 256'h1399bdbc46c439248a5dcbf9fcb8571d09487fa4c1fa1219ef97ed440b511d31;
defparam bigblockE.INIT_06 = 256'h807a1c586b465d0f0e4c05229b571ca22f8ac9875a5a038ffd007074fffb30de;
defparam bigblockE.INIT_07 = 256'h4dadc5aae41d57704d4739241004bda8dbe777ad5c08a4f62a208a485c908aed;
defparam bigblockE.INIT_08 = 256'h56c90fe1104ef61002e2100000645c62f0a1e544ee1c3144bb411a4bd8d34c93;
defparam bigblockE.INIT_09 = 256'h837e5a99df6e1393ff40ac2c55aec86776146874c9864e6fb0c71de2761ae263;
defparam bigblockE.INIT_0A = 256'h89f7fa2aa61bbb3616206fe851bbf6a1e654e07e596190bfaf15b22efdbeccbf;
defparam bigblockE.INIT_0B = 256'ha3349548c281e0ea6e1e931b02090d78ab7b6dc29226f674fd8fa805e15e67a4;
defparam bigblockE.INIT_0C = 256'h240045282a7c91e382f2b09a83047c234163b2c49e2a2b8e5f316c661a971ad0;
defparam bigblockE.INIT_0D = 256'h7feb8f1dff997c6f345fa7b255b9477b3d4807de990688acb86000b004b04000;
defparam bigblockE.INIT_0E = 256'h30d65f1ac235287ae621866e3628fad91707dfdae6492fb80ba30cfd86a7f68d;
defparam bigblockE.INIT_0F = 256'h74fffb72d2ff0c817af837746f793a5fb4e80a1ee6ab51d3764a81c91df9a2fe;
defparam bigblockE.INIT_10 = 256'he0e2960c2d1c800b71a0462521684df9230e4705e29b201e883dda393b438003;
defparam bigblockE.INIT_11 = 256'hc374190f4b7f08d6f36b567870cc34f96b2b094c21c5ba0a1b7f0cc9ef41b4b1;
defparam bigblockE.INIT_12 = 256'h55bf705ae4afedf1613a322d802340302100de59981d75614d6d9fb9f7389687;
defparam bigblockE.INIT_13 = 256'h6d16e50ce0a467308b487b8c369b685e931ff2f2655c7de23c1444172acb414b;
defparam bigblockE.INIT_14 = 256'hf804eff6fe33c82a8bb2affd0b7f7ff3441c5946116bad0e59b5a1a06933734a;
defparam bigblockE.INIT_15 = 256'hf19adad652ee8edbd219ee5d2eba79e5402cec99fb408db8a6637ffc9a72e1b6;
defparam bigblockE.INIT_16 = 256'h1281292294460925bb746ae1158ecb580d11d8cd090da016b1306abca156cdf8;
defparam bigblockE.INIT_17 = 256'h81827d00c4d093cf847837e321055cf38f4806321a1f2ae6f971b068b0c852e2;
defparam bigblockE.INIT_18 = 256'ha8dc3b1b884d73ac12939420fb4761faab054b8a37cff5eed8c148bfe1d3b1bc;
defparam bigblockE.INIT_19 = 256'h5b39fd43800274fffb723dff90276862f992ef6fdf49a29466f7fb95e55bb2b7;
defparam bigblockE.INIT_1A = 256'he8d1db4c0028215061aa6d8cad92f720462c236d0c19024e6725449ba82d863d;
defparam bigblockE.INIT_1B = 256'h0e5b7baeb2f9d83e40ca741f52c76db94e3e4e956b0f930c17f38f6af074a83c;
defparam bigblockE.INIT_1C = 256'h2767a053ea2c10e008b31166a29584c817911a820acd144001843e42aa7ce0c8;
defparam bigblockE.INIT_1D = 256'ha79b197dda70475bea0f4bde4551c744854f176c2795cd3e369245ae71cf9aa1;
defparam bigblockE.INIT_1E = 256'h294f3461e5bb2c9e6a5251c7edd3fe8c1f2ddfd7bf518d164ae653cd45f16177;
defparam bigblockE.INIT_1F = 256'h9a6fa4a09188fa56991ce475117d39de3f0b0b1c8e8537ff9c8e0810fffcffff;
defparam bigblockE.INIT_20 = 256'h15eab492c1b84906b925030a4000791247fb00b12f4fb28bf281e695aa03a546;
defparam bigblockE.INIT_21 = 256'ha834f6dfd907d76b16f4b54622c5ff029343929571d62bf896326d0d7a643268;
defparam bigblockE.INIT_22 = 256'hc630717c88adf421c3c495642c71cd348c7180926f635935330b91919263ee6b;
defparam bigblockE.INIT_23 = 256'h851b9032e93c5a39b63e000274fefb72daffb7efafdace20b1e972cc5b4f6b3d;
defparam bigblockE.INIT_24 = 256'h2ef32c6435bc92278e6d4577995ab12a6d0cb192f6c066200f680bad4bc24324;
defparam bigblockE.INIT_25 = 256'h1080f03fd1361247aba5ae2fbba8ef89838ce62459943fd81b8d69c9827281c2;
defparam bigblockE.INIT_26 = 256'h1ac118a5519a27a955c65db64b29c789d27258f48e8b10cdf42e9c1f0005b100;
defparam bigblockE.INIT_27 = 256'h8cfcc3657e31d974c351bde0fea20f0d52fde177ec33b2a3ffbacf555d09ca72;
defparam bigblockE.INIT_28 = 256'h8ede0422459136a55ef206b58c45b6ee5a8a7f76460a25a8112ae59e4c6eeb0f;
defparam bigblockE.INIT_29 = 256'h0c56a5e19f4ca2a16185eb6a37311b6b2a490801f5c0d63bd632d0bc49b6f8ed;
defparam bigblockE.INIT_2A = 256'hd5bbdcfced5db552ed08bcfaa1ec000096c900046610a4d3bf807e8631f7c9f8;
defparam bigblockE.INIT_2B = 256'h9375a357a1b1086056cfe2152bda5042881b254dd172bde1e5cfe1dd935531d2;
defparam bigblockE.INIT_2C = 256'hebe8098cd37b70ba3b50169b3af11f55032f0f5051ad1a4cb140f1fa8bf13308;
defparam bigblockE.INIT_2D = 256'h4ddda8a66718c4bbf82d2639db39ee4d800274fffb7000ff509332fa0d1a31fd;
defparam bigblockE.INIT_2E = 256'h908a50e586c552c988987fdb6627722ff6c0d0556119ed8c6a8a0fe064ad376c;
defparam bigblockE.INIT_2F = 256'h0e27000080c0c80cadb0d21e13692aadfcb5a618daf42052a4cc2490e3457638;
defparam bigblockE.INIT_30 = 256'hbb91026fde2140e298f9b022966a0c907e436508a3fceae3e181b231ea46ad82;
defparam bigblockE.INIT_31 = 256'hab41938fe1b3760965ddac9338533653961430ff979093ed4c3f213819c20ef2;
defparam bigblockE.INIT_32 = 256'h8fbbe8a59bbcbd092bea5edf162bd749a37eafbec54b742c87dba6c82e6c2241;
defparam bigblockE.INIT_33 = 256'h8c21a385863dad9589b98d2327ec1e456891416324ab36af249280109a9f1473;
defparam bigblockE.INIT_34 = 256'h933011bc8e12eb78790da960e6834fc93d1a8e96043d000000014412d1c72327;
defparam bigblockE.INIT_35 = 256'hffaa53a512bdd8566a325fa133223484f8e708e5ddbdc0eb86b295f5f94c611e;
defparam bigblockE.INIT_36 = 256'h3aaebfe63689274dabf9d0663e9bc287fedf64aacc1b9cb680df34b743e6048b;
defparam bigblockE.INIT_37 = 256'ha871a4f46da7f121764d2466bb6a1f822e3a398b4cdb0362ff807274fffbbd5b;
defparam bigblockE.INIT_38 = 256'h98c00985b0f68ac86cea3923022e000003b527795914bd53ffff0c699c138aad;
defparam bigblockE.INIT_39 = 256'h2c36a29c510a0f10000200001f8089a3147fe89c7722df76823f25bbc3b06bb5;
defparam bigblockE.INIT_3A = 256'h77463e70def7b5a2ff9a7ea44c2eb3531d7256d3940d70a2424952a7a7233122;
defparam bigblockE.INIT_3B = 256'h2856cd4af5b384b007594772cc03355a4c4f702be29e1352cab35e389b1f66a4;
defparam bigblockE.INIT_3C = 256'hfe0cffffffff67ff66729e17bfc76a5b7227e6fad9471ceff5648927ad104d8d;
defparam bigblockE.INIT_3D = 256'h60127d88946d674fa52cca7899b934901018fdae1b5a668741d40acada439248;
defparam bigblockE.INIT_3E = 256'hfe7056ed161d016962aac462a7e355c58901512c158235c7a979003b0000d003;
defparam bigblockE.INIT_3F = 256'hb16275f5dd1ced757d0878c3a65773f8f4ba6c29bfd45669fd8fb68152d2a86c;
defparam bigblockF.INIT_00 = 256'h7274fffb77d241324cb931a61c3f5ccb977e8584ab2859c8801ca7c474cd739b;
defparam bigblockF.INIT_01 = 256'ha54028908aede88c2cf86946ed73a00c2422cb4720626c5831884cda0349fe80;
defparam bigblockF.INIT_02 = 256'h92c28c87f51491c38e990f90132cdd259248d64ceb197f2990f14bee7a8f3adb;
defparam bigblockF.INIT_03 = 256'h0582d38485e9d6e227e91fae1f331da9083611040f1ccff8568234c5a6a8b5e4;
defparam bigblockF.INIT_04 = 256'h9a23525a770d6dc67262abd2331fa7ed3795f5e46a4151d6958e87f68f18bcd8;
defparam bigblockF.INIT_05 = 256'hffe9df675f4e7fea7a4766a3ef42e72da844ecfc994c1b3d8395fcfdd421e88b;
defparam bigblockF.INIT_06 = 256'hc558444e0f0b86130bcfa80b014434340e99752836dc010afffeffffffffffff;
defparam bigblockF.INIT_07 = 256'hc000a82043d071f7e0e473ad4e12c9bd09e7825d6c7ad0f10f4031226ac3f4ef;
defparam bigblockF.INIT_08 = 256'h3c4f1b4b92086bb509c9183f61748e1790ccd1820148e27f52f017478bd7871b;
defparam bigblockF.INIT_09 = 256'h37bb688315714567784f448053a9bbad88c7bbfb9dc967414e9e375d0a05fe98;
defparam bigblockF.INIT_0A = 256'h47d9035fff807274fffb0a36d001c7a35b3cce35437fdfd1daec15bfb2c9147f;
defparam bigblockF.INIT_0B = 256'h10ca2286dc29a030cc148aece0803d4f6726150d1c0d0d28cb3321625628b98d;
defparam bigblockF.INIT_0C = 256'h0cd5d46088a6945a18197ba31fa01a7bab02949b88312c664a1a0fda49088076;
defparam bigblockF.INIT_0D = 256'h06a153776d7a8141728a625a472309672c3d8446005118084068f6933239b738;
defparam bigblockF.INIT_0E = 256'h308477620b567348aad9b6317a54804fa0cc10af7f674030aaacb1d6e72d82c3;
defparam bigblockF.INIT_0F = 256'hfcbfef6f3b6ee6eae92a95db3ce0cef4c443ac044b9a413757ce79afe540cd26;
defparam bigblockF.INIT_10 = 256'hcdb818a6ed8828d252652648fa4fdd4740bb0cc141e4dfb44e3600010000a5a8;
defparam bigblockF.INIT_11 = 256'hb2ff6bcb80560925820065a70947407e5ecb6224a838657871caab813eac9890;
defparam bigblockF.INIT_12 = 256'ha1f085d2ea9a36d4414d91688b4cc9f515ad35375bace1e73ccd1cf2d0c90211;
defparam bigblockF.INIT_13 = 256'h9ff9ffa83d871325a670677b3d7980f1e134ff99da7dffcb27e33217f4bc14b6;
defparam bigblockF.INIT_14 = 256'h34c53c4011eb43d902d7ff807274fffb00044c00007af4e8dfed8b3f2b99bfd0;
defparam bigblockF.INIT_15 = 256'hd05fd7cc975d3c0a6eb2071baa298c9293ec40c025b16466c90fa00a24271b23;
defparam bigblockF.INIT_16 = 256'h009950e08f0a34de3dff0987d769c290f7624da9a8a7a66ee10e81c3c8eb42fd;
defparam bigblockF.INIT_17 = 256'ha1880cd538cbdba0d42d8f0356254647e08a020eb18d01e8804010009130eb45;
defparam bigblockF.INIT_18 = 256'h6a57989634c94fa536b59a93e271be8ac6c5659526094c2b01343e7b168ce7ac;
defparam bigblockF.INIT_19 = 256'hf7f897f4e9479b3aa9ababd800447729645f40a6b3b08524796d1ef5a04a1dfc;
defparam bigblockF.INIT_1A = 256'h36a8a8c35294aca99890934a2a46fa08ffff51ff06cf656ac2ae1f7eae71edec;
defparam bigblockF.INIT_1B = 256'h1894d9dc0310203d00002004846be8884097b5b6a626622c0e4836668eb6af76;
defparam bigblockF.INIT_1C = 256'he9890f3dcc5426774efa06e0ed5a4b9f4dbbad48074cc08f0e57a6796407a76b;
defparam bigblockF.INIT_1D = 256'h5ce66fa987e690d1bcadaab233e0eec584f89b95ffa9ac5aa558ace8b2969cb7;
defparam bigblockF.INIT_1E = 256'h7c4a24ad9b3d34c43db0d18a3e5902ceff807074fffb3f82ed7982b7a6b706cc;
defparam bigblockF.INIT_1F = 256'h35d69fdf01201722caa59ef70e0f5e55ab85a1f1e8c313ec80cba4516747d8f9;
defparam bigblockF.INIT_20 = 256'hbbfc0054000087aa07fa22430a2b8e3f755a4a508b2a7615189024095d8e447c;
defparam bigblockF.INIT_21 = 256'ha285b30355ab36341a7055eeb26865a5c374368974ea14ae131df408f9785184;
defparam bigblockF.INIT_22 = 256'h35f6281ab1181442a410ed55a3639607c4d9088269b7515a197893d8ea5e526c;
defparam bigblockF.INIT_23 = 256'h29ff09c23e860a969166b21e7dc790ee0afe7fc8ebabe4650ed4c5628e2cc590;
defparam bigblockF.INIT_24 = 256'h180e502cf48203dc322a18ae5d166a7cd066d43038c11f85e6aa0002f800ffff;
defparam bigblockF.INIT_25 = 256'h49185c4501042789a446476cdab60a95000000007283c999d3fd88750cb1912e;
defparam bigblockF.INIT_26 = 256'hd3bbc3c548601fb52f981f36075220b27ea1c3cf01f841ef1b0691780129fcbb;
defparam bigblockF.INIT_27 = 256'h1517cb7bfc66fffffff8ae1b858b6f8a6fadcebd7ea68effefb421b8ae2aa4cc;
defparam bigblockF.INIT_28 = 256'h51e0e7a40d640c65a982273022bbd824e914d9516d4d000374fefb72aeff1e6f;
defparam bigblockF.INIT_29 = 256'h1d4bc40c6efaaaa063a1893bae9b003fc2b0e585c1c320390896928eec88788a;
defparam bigblockF.INIT_2A = 256'h26e1ae5d809c000000000100499aaa00c277b352aa9365842616c40412048bde;
defparam bigblockF.INIT_2B = 256'h2b0be0b650c3b92242c83e0a91312dc6c294c12f4637d063a2b85f098e40bf55;
defparam bigblockF.INIT_2C = 256'hbfdbef1f8f129ad25f2f5db9fada9d5c053a6b1d41784fb299087172466442e8;
defparam bigblockF.INIT_2D = 256'h3ae5d38bce75a6d8b93e66637175588ff98d3ad2ceb245619aa9323ce44e1e5a;
defparam bigblockF.INIT_2E = 256'hfffd1fe37cef1ffcf5ff0c988d8c336c55c5a45ffbb19e9e5abbff9c62f3718d;
defparam bigblockF.INIT_2F = 256'hffff81ff70cf3e26f713f4bdffffff5ff3ffebffadef358fa7c6677af37aa969;
defparam bigblockF.INIT_30 = 256'h1231c2330f2385a97a8c5da11540561268627f3cc98a2187ecbda285dd22fbf2;
defparam bigblockF.INIT_31 = 256'hfb7278ffdb343b528af23f674d9ab138903015ccc6d131b492ab246962f37595;
defparam bigblockF.INIT_32 = 256'h98606c1a9288000054c40d610c05c9740930c2bb6828862c58194443800354ff;
defparam bigblockF.INIT_33 = 256'hbc1ae63c005ff52c6bad148f6687976dd6ed39e5e090213445500ab3000c01c0;
defparam bigblockF.INIT_34 = 256'h3295fb5a14cd7769381ddfccf3ba37cf48e0de362e4998a2707539a8a2806ac3;
defparam bigblockF.INIT_35 = 256'hc0575295a14c82c2695342202f90f401da6cff730ecaa1bd926557d2c5208cfe;
defparam bigblockF.INIT_36 = 256'h4a3cfbbc9656b706154a8ac50820bf90cd05390b1bb11c0a94457333e3a4e96a;
defparam bigblockF.INIT_37 = 256'h1572d07ce636fbb2f88e14551de5e3f98f6f6ca6d2b923145248f18c471ded31;
defparam bigblockF.INIT_38 = 256'he11d8caadd1593ddb12dbbbb05bff4aa6a86fa7886dd5a5bbb3bd35d1591dc0b;
defparam bigblockF.INIT_39 = 256'hc7682fd2ffc28d7fa7a12927afc2eee5ffce977fa1a46e0331974b25578d97cf;
defparam bigblockF.INIT_3A = 256'h402a1442280fc24c3f8abb525538ccaae500d32afff9ffff90014de90cfce54e;
defparam bigblockF.INIT_3B = 256'h4164800574fffb72afff8386258852604a5c413c08bc2e3a8a9ae0ef98023f2d;
defparam bigblockF.INIT_3C = 256'he22d019900121ec02b8b078f0001399c915c1cb9bc00e2c743ca00413de05736;
defparam bigblockF.INIT_3D = 256'h0919f7ac19660634d2852720015c925212224204e13a194b62b250cd0a042c8d;
defparam bigblockF.INIT_3E = 256'he1e62eb841e3977b4270ec725235411d8ed4810b5b9a87c8300750ea108aa056;
defparam bigblockF.INIT_3F = 256'h79976dc863d6e356fddf7d75553277cd577c476f70dc7dd7495518646bfb20f4;
defparam bigblock10.INIT_00 = 256'h46f92492a6b7bc0070c5e9adc045fe13e63d2e78dc9fab32cc4c0f1775c78ebc;
defparam bigblock10.INIT_01 = 256'hb05ba6d0bbd8c51db7aee84200c2748005fd6846520aa910a25893525b68f252;
defparam bigblock10.INIT_02 = 256'h4d315253ecee1ce29462978f25f0571269b4f2dd9cb7e044d5635a7dfbd9ca15;
defparam bigblock10.INIT_03 = 256'h0f5a19f5ab33e6eb7ed7367e00f731ef5db32291bcd330cde2c16e2d8ab34001;
defparam bigblock10.INIT_04 = 256'h4f3efc12a4a61b6d85134c02f59e7e57f31d5d178b1a1b2d4d5550bb2e2ef7ff;
defparam bigblock10.INIT_05 = 256'h0a153d00dde75e5000037482fb7052ff171b00154ac027236800b0930ce9abe4;
defparam bigblock10.INIT_06 = 256'h3bbae443ca5b6aa5ad5908bf008c6ee84905d8e8260c25770cdd8c00bae0221b;
defparam bigblock10.INIT_07 = 256'h878786853239e466da0cdcb1420c645dae826ed14e3e54ac5084f2bb2cb596b3;
defparam bigblock10.INIT_08 = 256'hb420223c98f5eb1f34c33b79e7b697b48569b3b9d50c85fdca88b9be46b028ad;
defparam bigblock10.INIT_09 = 256'ha32f5088d9ed7d00db4a51b6a491003047489dfe9aaa9953ee7b25a339b41801;
defparam bigblock10.INIT_0A = 256'h686a8edb1124f52a7980e236a3a9b5679c0e0a92711006860e479e80b4784337;
defparam bigblock10.INIT_0B = 256'h5d5adc6a311669bef3b663320597bbd04a6c3528f645e392106e588ba87e1db4;
defparam bigblock10.INIT_0C = 256'h4b1db3a1851730d4ab14fcdcec3c1f5ef3769e1cfa7522f3e71796756f24a564;
defparam bigblock10.INIT_0D = 256'h1e263a304f3ed43b1132c9ac7f26d2417236486302559ab6826cdf336ac3fb19;
defparam bigblock10.INIT_0E = 256'h9da1575f9ec6e85da9b926090ae83b14ccd5c376d09439e8000949a0326a1640;
defparam bigblock10.INIT_0F = 256'h000c00221bbd15021dbae185455d03278f807274fffb9bb33ec219e8efd18494;
defparam bigblock10.INIT_10 = 256'h526a6630974a4a3678ad5a8a4a11364138590d80f413086ec85e147877e69535;
defparam bigblock10.INIT_11 = 256'he5fcbdbec77763280d74ad9d6e0e84b674a16a93332e2b65ae74a7e1936a32d5;
defparam bigblock10.INIT_12 = 256'h5880a800c006852b1f42944a2c0e6e0523941b6d1049011c5997b2facc611ecf;
defparam bigblock10.INIT_13 = 256'hd4419fc9ff88c0f7b89e52bace7c90ffa073901fd0be3d50865c8ab8a89c070b;
defparam bigblock10.INIT_14 = 256'h94d67d4555c30cd4d44f1fcac3b6e07c3b3d534b3bf94afe22d9676f82bce9bf;
defparam bigblock10.INIT_15 = 256'h0c28e82a5bfb4d9b85c0ed7917512db60c47baa307d8f72a55189a470447294a;
defparam bigblock10.INIT_16 = 256'h9c6d20226d860541293a49e60611e78450b6a463236d2949010950094e1b7040;
defparam bigblock10.INIT_17 = 256'hb728798223b15f919d3a2ac9c2b57c14f5384e0c4d31ac09cb5d116a0019a000;
defparam bigblock10.INIT_18 = 256'h51e3a29d63149c81acda9a078cab50c109ea53d1c5119e3d8e06bd984c6017d0;
defparam bigblock10.INIT_19 = 256'h24b671864d19180d00261b8a124115a269874cdc03189f807274fffb13b4cef9;
defparam bigblock10.INIT_1A = 256'hf6d733bb0f95a2e9f341d16cdcdfb5225b617a2a99d5f35d88203400896ee05d;
defparam bigblock10.INIT_1B = 256'h9cc18bf777f000bddc3f0e114e189fa48e3619241b61e00366644ae7da1480fc;
defparam bigblock10.INIT_1C = 256'h2b356cf69fa1044a8a81547ab51960f09eb05a14b92680125380c1b84e00cdec;
defparam bigblock10.INIT_1D = 256'h1d2bb4970c6e6d67a056f04f4514ed0c6aa16e198b0d0f859d0375682148dbaa;
defparam bigblock10.INIT_1E = 256'h19813c792cf86b59dc1050e3c3406ca96df02a3f04ab2b693ab16a8bb34d76fb;
defparam bigblock10.INIT_1F = 256'h014b94005c540a01195fbc6b3df787fd6f6e71f5295f20c26da94924c859a801;
defparam bigblock10.INIT_20 = 256'hca98de93e384f7d2dd09a88bc87680c73fc4d1c4816e86c12176440d32a45981;
defparam bigblock10.INIT_21 = 256'hc6759b3b3da97fec83a63d386516c83a5e5d9c295c282adefe06f4f6be1fe21d;
defparam bigblock10.INIT_22 = 256'hfffb0104f81844a9b241d43b67088e160739f4b36da876a64f31d2d5517f35f9;
defparam bigblock10.INIT_23 = 256'h2801096e00609c5671a4c4d90a0b00685b8d1a82155a69874a5c0343af007274;
defparam bigblock10.INIT_24 = 256'hca1456e22ad37327eeb8e0d911b56d1df4223c13324a836745066d6ba31b1848;
defparam bigblock10.INIT_25 = 256'he7dcd4e01e55ef50068b0fefbac99281feeecdb0f192c0905c60028500000220;
defparam bigblock10.INIT_26 = 256'h3ff9658f6e3c3ec3b761e271407ef8d61cad6ff02c59e29ac51fe384bad50202;
defparam bigblock10.INIT_27 = 256'ha2e0bb415d62604d614e78ee9672ace94dac57e38ed4eeb93cece7df088e8569;
defparam bigblock10.INIT_28 = 256'h9d3b1deecc632669054c020014b08d55c78f1fc541298471b45ddc8d00482040;
defparam bigblock10.INIT_29 = 256'h57abfdb8bb918339519e97b10d7dea87897f95fed08e6bd61c5c506d37c5a4d9;
defparam bigblock10.INIT_2A = 256'h8ab90ee465904815f6f9efd02b21019c5851405df50528adf63c001ac6cc6926;
defparam bigblock10.INIT_2B = 256'h105dbe03b6262ee978f746842465e48d08b81404d4605da5cacc2357e24f2a2a;
defparam bigblock10.INIT_2C = 256'h030dbd807074fffb78581dea8a66af3128368c4518a3f2d5c2f9005609402ca2;
defparam bigblock10.INIT_2D = 256'h29ee9ea38c003400852ee046a051714411352c0c04623b8a2044436850c942dc;
defparam bigblock10.INIT_2E = 256'h8f258850c3a163175491fe20f1525233d1950d2ca26990f226abcd118f09fc3e;
defparam bigblock10.INIT_2F = 256'h91d544b399c855f5b436a0d972ada54166ec7a96bd6f0872704cdbe6c32c5cc6;
defparam bigblock10.INIT_30 = 256'hcddd00271432112bd005a1316915b8db806961421e014f17a8c2dde872e53edf;
defparam bigblock10.INIT_31 = 256'hc9330452cb2a94d308904a2b002548025400c2000a44e452b1743f5041ee0590;
defparam bigblock10.INIT_32 = 256'h471530b5a77f8d8f2e3e1fe6c033e16c8c23ad4e87b96ea59b1536684a6fad36;
defparam bigblock10.INIT_33 = 256'h0b78c895810ce500a4cfa247bd060a11561f2a4219bfaa8047fc2e37ea1f1a4e;
defparam bigblock10.INIT_34 = 256'h161f815d5fb11a6992370002c03c0519a32a8a1fba0764474cc40605d9461a90;
defparam bigblock10.INIT_35 = 256'h30a78bab32ad8fc6211c4e3db05838b02990400101a448452c80ab18e940b6c2;
defparam bigblock10.INIT_36 = 256'h081225175cd1d33e000274cefb722aff80b96d5aa8bb077dd2ebe39ee6222c6b;
defparam bigblock10.INIT_37 = 256'hf1d83cd194cc8b80f30631f60194ee74888c51e0a62075734d19490c9d00c16b;
defparam bigblock10.INIT_38 = 256'h32b3846f31ce1cd4e933455aa2189c63fd67b320733fc1246182883f453045d3;
defparam bigblock10.INIT_39 = 256'h9d0ce77a692426db112ea70322a819c607e5322953fb6391d9aa636d7b4c57b2;
defparam bigblock10.INIT_3A = 256'h5a98fbdb4c8f95637137e08a9dd1496901431200000a240f9e612b24e935a0f9;
defparam bigblock10.INIT_3B = 256'h1725cf5f48440ba6ffec2b6684a7d7af14b6db1e5c48bc7d19665ef058cbfdd4;
defparam bigblock10.INIT_3C = 256'hfe15c49f4eea67b79482bb8991c1f7a99802ef504d77edb83065e35e98c9aee8;
defparam bigblock10.INIT_3D = 256'hb68b148d0040bc38e982b243ca84af047ff8d78cf05d865a8a49f8bf8dff6ffe;
defparam bigblock10.INIT_3E = 256'h97104020c0483c1e0f036b8c844750f3d62b3de98f43d0a6adfad62549330b2d;
defparam bigblock10.INIT_3F = 256'h32b7f0ab6ac7b4287a5d26e2ee333d51433476b5a5fd69931ee82e1bd3388648;
defparam bigblock11.INIT_00 = 256'hc5307d0c21abd0158b1cdbe92a33000374ddfb72adff600dc774d9d4b246e367;
defparam bigblock11.INIT_01 = 256'h6fad37f462865ffb4234ae9a6727bf5da8271494ade85006b608a62c6d6f0d35;
defparam bigblock11.INIT_02 = 256'h4200558975bddd5dbff5295ab3fe5b41aad2f7fe5319fd6ff8d7dd8fa2f91d0b;
defparam bigblock11.INIT_03 = 256'hac3448b9d17b00200020004092896c213154fe7d02f5bb0a9843ffd202773200;
defparam bigblock11.INIT_04 = 256'h53e7cea652b3d971d4e0be1d61dca235d2a8449ca95666b49cf10891cc242e96;
defparam bigblock11.INIT_05 = 256'he54fc107ee5ac95f2049c8ef1d45fa72301fe9d7aba9cf013745efdc0489b69f;
defparam bigblock11.INIT_06 = 256'ha7b199d35ad472a385852d5ce9a3b6aaac8e335ddfd43a908f59b6ea17fad8d4;
defparam bigblock11.INIT_07 = 256'h7e14a21383379ae459be425384a99a89ba05927449260b1340007c04aea2746e;
defparam bigblock11.INIT_08 = 256'hfb33b6a2e9154a9cfbaa959ecaa9aa10c61e4520fe4cb3dc4bda00040000d802;
defparam bigblock11.INIT_09 = 256'h98d54a48296b4d74b110d950318b877ef397ad71ce3c65c1311769acda92545c;
defparam bigblock11.INIT_0A = 256'h47a0f9670c48251e3a0502bb2220e92ed9d17e33000374ecfb7201ffe425b75f;
defparam bigblock11.INIT_0B = 256'h84f52fff8f9e5afff8e7e36f56ea2cc506e6b88ad6aa9023160c6cf05406b888;
defparam bigblock11.INIT_0C = 256'h846edb608f506ab10a750201c915b7d96a88b4b7170c194e5e6aa88beacefe5e;
defparam bigblock11.INIT_0D = 256'h218f59528d25246bc16588f518b800000000c00002001c07a360c6525eaa0feb;
defparam bigblock11.INIT_0E = 256'ha2c87189d7d6926862d362b944bd57b771b0f1734d9ae1e36da61b6c89445d66;
defparam bigblock11.INIT_0F = 256'hf2fa020e846a5afbb9937e2b61b3c288d4540f3c851a37ba7b6e2facf6324cf5;
defparam bigblock11.INIT_10 = 256'h5557000d0d00a3f015cb6998e080b6f987010b5a61a5659627712b6a5f443a97;
defparam bigblock11.INIT_11 = 256'ha4f116cf32db02ab0000008005088ba8540e0517f3e62f7106936289c3142492;
defparam bigblock11.INIT_12 = 256'h4cf50966aadbaf1e1e3da4884c7ff97f82b61ba1149b8523914b07ea41402e5b;
defparam bigblock11.INIT_13 = 256'h0aff59339f5c723760f5902c462ace3e9c82baa371931a87faa1723acbe03f30;
defparam bigblock11.INIT_14 = 256'h6be45c050b808c3d255f0dede908fd05e1aa301beb1657e1865e800374f3fb70;
defparam bigblock11.INIT_15 = 256'h5efbbc16f8629dfcfbff054fa8b93cb176a13647bf09925ff27f57c399e565b0;
defparam bigblock11.INIT_16 = 256'h068700002000dcbaa42d10de7a4c0685cc9362ee10d5a0ccbaa800aea000e100;
defparam bigblock11.INIT_17 = 256'h89750623bc54fa85e50f3c53d31b7198304755a1595d68fe050dd2e1f1c1ebe3;
defparam bigblock11.INIT_18 = 256'h57344c91f62fa1fc0c7a85473ab243162767ad5db6d25f74e687ac89d11a0283;
defparam bigblock11.INIT_19 = 256'hb2366ea7c2567001e5b12353e21e022a2a5d40b09d978b81b8f956672ee28162;
defparam bigblock11.INIT_1A = 256'h9b68efcd93a23b0233bb0430814ba0a42aae555f0015fe00ffff88ff60f3e38e;
defparam bigblock11.INIT_1B = 256'h97bdd76b17506e92dedac1bcedae4ecc69e2b7ae1a90a32ba7302ab000001c00;
defparam bigblock11.INIT_1C = 256'h032ea69973b75afdbf34ac7352ade2a63372b87df0c10b65305dfa8d888034c0;
defparam bigblock11.INIT_1D = 256'h0374f4807274fffb721b2a370a6baf354f652f9d532ba6153c15cbae9142d3eb;
defparam bigblock11.INIT_1E = 256'h2f88f5729888303786ace863b0ab61a76cc9160d05e67b0c184116a869e843d8;
defparam bigblock11.INIT_1F = 256'h7f18a06ad3001d47c5860e484db5b513000121a024797318481d57fe332f93f1;
defparam bigblock11.INIT_20 = 256'h7b5298ea93c4930342cbdfc6602590993c1550dc0000db00ad77b10f945e586e;
defparam bigblock11.INIT_21 = 256'hbca112328a208bc959a112699128a362f939e9607522d10b779cbbbe4d7c2989;
defparam bigblock11.INIT_22 = 256'h3abc8e6a472c0f7607f62c914c5106b0b431e42d64830e3cb7cfd649ca661417;
defparam bigblock11.INIT_23 = 256'hfeaa000bff01ffffffff3e8f6d4389c0c9b90a2dd097194a7a0e141b56fd16d5;
defparam bigblock11.INIT_24 = 256'h2843984d91b3006000002e344504457b78c0a142c66d60bf164261e98b0f84d0;
defparam bigblock11.INIT_25 = 256'h281d142801f88f027119f28e430366881708c3b0420fe4992cce85a0b98e21c4;
defparam bigblock11.INIT_26 = 256'h5472d69580bce8e2e435ad74db089195c93c90f8a03c3a22e2ac41908c090ba4;
defparam bigblock11.INIT_27 = 256'h42f839ec34d70377fa007274fffb78ff6e3dabee857f29f995fda2cae5260e3c;
defparam bigblock11.INIT_28 = 256'ha451f0356746e5a8bfffb0c8a86786abe06eb0af5c671127320d1969aae91801;
defparam bigblock11.INIT_29 = 256'h8b0d4f4348ef4b628d3f75587484d2dfbecab9a88a49322400009000d2ec5fe3;
defparam bigblock11.INIT_2A = 256'h3f8695567e2b59228fa5d7436758994c6c41615b6247042408000000bc04a71a;
defparam bigblock11.INIT_2B = 256'h0e3efdb7da36ef8d5e90ad7b46dfd5a44df73b790aa8d79bf597a6e6a531bb5d;
defparam bigblock11.INIT_2C = 256'h6ffb8c7b2ff31f1156c9be257a3f1b8bb7ffee14111e6397c9314dc6723427b2;
defparam bigblock11.INIT_2D = 256'h0bbb4fe17aed2e5063deff5de77f6a67fff7d7ffdff79b75d2f6bbfba7d6df54;
defparam bigblock11.INIT_2E = 256'ha042085a4b1d797910b5b09d6cc339d0c272233829575478a555c0aa4abfcdb4;
defparam bigblock11.INIT_2F = 256'h54a378442583a39158e385729944ce0710f34a2c89a00190884750ca08a07331;
defparam bigblock11.INIT_30 = 256'h716d058ea1e3c30453880ca69954c42c1672c6f227d20b48cb83343487214489;
defparam bigblock11.INIT_31 = 256'h0d2caad91ae115b899e945d60390ff807274fffbfce64e54f3499c8b697d0b34;
defparam bigblock11.INIT_32 = 256'hfd693e6495cdd42bcc53b3babe76baab6000769e86ab2079f4005a74590f040d;
defparam bigblock11.INIT_33 = 256'h9e547128d47c4d84a5ab16f22a16b85ac51313d26784970abfa00d21b2c95f57;
defparam bigblock11.INIT_34 = 256'h5c81542f9f30b6345a1394fbedada8a6ce1e0b278eceda77c1f7a8bc4978beae;
defparam bigblock11.INIT_35 = 256'h12712e4216a3427118e69c6e166355552aa919d0439bdffeab71ffb37ef79d3d;
defparam bigblock11.INIT_36 = 256'h17d5e832a88a2c854e9188d963fa200cd07342d146253c0e213e428e5d9d0620;
defparam bigblock11.INIT_37 = 256'h8ea46f86f3610000534c00c038c3b2ac1e5fa4465a8d3c98e7d32ad350854a41;
defparam bigblock11.INIT_38 = 256'hde0a6711c5518f97072258e124311d428f23340837521fdf1e925116c8909d2a;
defparam bigblock11.INIT_39 = 256'hb3fcf1b6eb8fb97b6d7f78e26620e6ee1bb8ef6b1491cd4f3067f86676ef10f9;
defparam bigblock11.INIT_3A = 256'h5354ffaac16baffd971f139ce3c65533936d36d6ff2da3fed2d049d5cc73cdc7;
defparam bigblock11.INIT_3B = 256'h5a18050f0011c7a4cad23d23e0009e3d4dd6040aff807054fffb4f345290ca74;
defparam bigblock11.INIT_3C = 256'h5fd903c4e47a0b3b5e3b4f27000084000b80b8bd7c52f0004b1e0f2b091af600;
defparam bigblock11.INIT_3D = 256'h9852bc9ee5f791df24c0bc84a1ffa786c9943825a7b6f47e07b2b0a9787c0865;
defparam bigblock11.INIT_3E = 256'h21a1a0847830dbbc3347dbc44e2e605708691031569806280d66d042fbec18d0;
defparam bigblock11.INIT_3F = 256'hd755000d36aca7170e3e2848ab98dd6083e1db10d506b024acffeeff3deeaed3;
defparam bigblock12.INIT_00 = 256'hd89799f70aa88e413c0a90257084125b1b9288414299b1cc209a42c952a71f27;
defparam bigblock12.INIT_01 = 256'h81960a399a88a838369d360a931c27c133da4c72d758477b8eab7b2f484d9ff1;
defparam bigblock12.INIT_02 = 256'h7f45ffb9b5975fc2b19e52fe217917ffdb920736867d52557ce3a9335bfaa15e;
defparam bigblock12.INIT_03 = 256'h9a4949c402dbf8311dc76066b28800c08b2009c3b8e92f7c919c6f1a2a5e7553;
defparam bigblock12.INIT_04 = 256'h56ffe2a856e0b50d503e29d30003cb0a13b5ddb0d2899d5c7809dbce39d92099;
defparam bigblock12.INIT_05 = 256'hada45085d060232c236d4d79000066e3812b081119005b672d56800354c3fb72;
defparam bigblock12.INIT_06 = 256'h3098c9b2696ab83b8bdf1e0bde7465e52d8c7bdfde87f1b08548b4ad8151608d;
defparam bigblock12.INIT_07 = 256'hf7776df36c99e9878fd841120fff523d631595e836995149d456a08c123b758a;
defparam bigblock12.INIT_08 = 256'hd9328a12f540862574a87ee774883eb2c9ac2522f62575815cde9d4ff3f35b76;
defparam bigblock12.INIT_09 = 256'hc5db3b09e5ba3cb08a3500397088a79a2901771db667f2c695d6dcd0491f371b;
defparam bigblock12.INIT_0A = 256'hdb706aaaaec521997fd62c18aff6fa924110548e46b89d5b1225ab3f12285006;
defparam bigblock12.INIT_0B = 256'hbab98f4e516e5918d95c9eccfa5275ac76311b7ee6b5626aca2fc42eb1828b6a;
defparam bigblock12.INIT_0C = 256'h1782c079d42a71b6451b5a29fc022fd9870eea358c9d9d5d969acd764a8a9edb;
defparam bigblock12.INIT_0D = 256'h1202b51107b1cadff14985c73937cba4b0fcd1890c2c6000438b8042f46a4109;
defparam bigblock12.INIT_0E = 256'h000374d3fb7257ff21fe88de11c2f894ff26896780df2604e0016bacbc5d2eed;
defparam bigblock12.INIT_0F = 256'ha69e00b31018aeb44f05d568879c05754d392602ad00e16b2214881ddd694d5f;
defparam bigblock12.INIT_10 = 256'h3ca1b58ef1c1fddbe5b1fc488ff71d93a7420d917eac82667624cecb94e9c06a;
defparam bigblock12.INIT_11 = 256'had66ed8444f6004f34b9d8581af772478284700819cdc5dc976373083dab1a57;
defparam bigblock12.INIT_12 = 256'hc9b7b3eb235d62cdb324d0c898b14a61b40095a5400a555e141a0c948a2efc9e;
defparam bigblock12.INIT_13 = 256'h377058450e34e624c71e59ee942868846615a694a9e98963331122563185a7c8;
defparam bigblock12.INIT_14 = 256'hbf25d4d3febb6a8ff08cb66fd884de4fcc44d57fe8a7a54f400c77e7562be1c7;
defparam bigblock12.INIT_15 = 256'h0e20be776c9685e1b50bfb6b2ddad90866b9eec95fff48954422838fd4969dec;
defparam bigblock12.INIT_16 = 256'h600fc32837b4bfea194bd203d95415903227e20351ec001898c073365bab2ace;
defparam bigblock12.INIT_17 = 256'h20fa5b10f0cf93d9cee00491a71fab6db255404cf06c8570acb29c44e3e09ab5;
defparam bigblock12.INIT_18 = 256'h862ddde11e5b000374e0fb7215ff7ec6a9ba02c2edd11a3ee0a1dd1031f91af9;
defparam bigblock12.INIT_19 = 256'h612ee37f1f576fce415f231e2ee87a0c7a60449817774c810300bd00c12b2a11;
defparam bigblock12.INIT_1A = 256'h3070d4ce2dfbc49d56629348b5631c6d2aa70223040363b30c1f6b7522e3c9e8;
defparam bigblock12.INIT_1B = 256'hc7373bc6fb0127b1d82c25d6240000198c52916aede2105df18d1b53d5b78016;
defparam bigblock12.INIT_1C = 256'h10ed89b4d8a41f38a298fb913886bd14647841147909302ddd63ee6f737284e0;
defparam bigblock12.INIT_1D = 256'hbfadd91fdf31a55868e6f9d476b75960f43db491839709c23698396efa2f72ac;
defparam bigblock12.INIT_1E = 256'h218c6ba5f3ce8db5049c4480101a172471e52a379d73010035ea35d57fea87d5;
defparam bigblock12.INIT_1F = 256'hc40e7a70472c048722002848b6683d6bbd15eadd1b48bef980a6b3e2586eddd0;
defparam bigblock12.INIT_20 = 256'h74c67cefe6b1ad0dbebe6d5b2c9afbde154aac6ceddb296b29566155c6072349;
defparam bigblock12.INIT_21 = 256'hf3bbbac656fe6f4063585ab07b5c27d585aeac7253158bd3d30ca96ab61c22c7;
defparam bigblock12.INIT_22 = 256'hb90982cb121c23165dd1df49000274effb7052ff9894a32a4377b554169a55ce;
defparam bigblock12.INIT_23 = 256'h4eb3d487dabf931aa7e24fe766c3100900a0eee88a8dbe20449c25774ca12390;
defparam bigblock12.INIT_24 = 256'h424d9a54c9f2853d1e315ae2a1906ecefb8a19c1372dd3596e83dfff8410bf88;
defparam bigblock12.INIT_25 = 256'h129786a9b039452df9bdc9ea13960698edc291a13af16116770e2859a04e4517;
defparam bigblock12.INIT_26 = 256'ha1bf5c95672218f11b3adffa9b5e20e9753c440a39c1ca49bd124f3dfd5a4b2a;
defparam bigblock12.INIT_27 = 256'hfffffffffffff57ffa9ddf2b4fa14c6eb72ffe56cb7f4115e3fd925e12c79180;
defparam bigblock12.INIT_28 = 256'h4d43a044cf3606133dfed67771b604008000ffffffffffffffffffffffffffff;
defparam bigblock12.INIT_29 = 256'h0ed18a1d7d278caaac35009f790808629eefa8805e1581d2841f6c0f7e69d3e6;
defparam bigblock12.INIT_2A = 256'h637f9b6e721c33bdca2e72eefb1ef55896cc2518d2f8f62ed2239b7c0b953e7c;
defparam bigblock12.INIT_2B = 256'ha9bc0a5ff485dbdfcd5b5c1b32eac4e99db7656d171df5bcac7df02486724252;
defparam bigblock12.INIT_2C = 256'h71265541640d18287b871ee32db0518848dc032ef9807274fffbfd1a2a68ca43;
defparam bigblock12.INIT_2D = 256'h1c1c61b62296bf39e46d4400ead44feb1bbf5bf429bd8cb918240ceea07f3cf3;
defparam bigblock12.INIT_2E = 256'h285a15400000802689005f96451abcab28f33847435ccad9fe0feb108fdfb82c;
defparam bigblock12.INIT_2F = 256'h121938cd6b25908a558a27e1e0153d83028b76496a300e36f34668a90f174814;
defparam bigblock12.INIT_30 = 256'h31186ccd2775a0f4fdc63291b67f812438eaa223bca4f3f7c0b9a6a58d57b150;
defparam bigblock12.INIT_31 = 256'h9fffbfe22d7e522c3d7495fa27db35558e86fab27d91232a634556cdaee5a0eb;
defparam bigblock12.INIT_32 = 256'he41069ed25880c722b149ef7c53513552caee45935a0dbee2e460088fffeffff;
defparam bigblock12.INIT_33 = 256'h1c02bd9aec30e29bda5c1599ba2feefa9588dafb0eba1d6484000505d47067c7;
defparam bigblock12.INIT_34 = 256'h4364ab11ecb1b9ba9bf87553deb19961f6edbd324a31719ddd3dac6c78e967d7;
defparam bigblock12.INIT_35 = 256'h5bf4542fbd59f433c70dcb6e91aaa063c3c03f76a531077676ccb216ba4c6147;
defparam bigblock12.INIT_36 = 256'h0ded00892c5e6a46b523824b19833b5a25031470898941da0361fd007274fffb;
defparam bigblock12.INIT_37 = 256'h3bd6b00b84572590608f7fb9c6db082512009630835faf6fdcb236f78e404c67;
defparam bigblock12.INIT_38 = 256'h2f590b4765b9de35e38e070940000820e95e950990d11d36fdba721155d0913a;
defparam bigblock12.INIT_39 = 256'hde4d92ae569bdb4f434fb73354cc735825a642d739f7d12ea366c7cd41be9611;
defparam bigblock12.INIT_3A = 256'h0dc2c7cb3b3144e704a8a00f47dcd6836d855e5b02e9d125998aa8a3cb676117;
defparam bigblock12.INIT_3B = 256'hff80ffffffff5039ab5c610537f284422da396ffd2f995ac4d29a5cef942afeb;
defparam bigblock12.INIT_3C = 256'h3a4538e6877c7f63a9af4bb02bf7f6a36ee4948103d22807b6b3fa986e461014;
defparam bigblock12.INIT_3D = 256'h6079ee3bba09ae7afc290b6c573d63540fcbee8ac12c5cb9946a490492c07fb8;
defparam bigblock12.INIT_3E = 256'hfb511d516e1ed9a5f6fff76be9e4b6c2e521dfceedfe78aaee998a18ecc455d4;
defparam bigblock12.INIT_3F = 256'hff807274fffb475d8770bc2a95d30a9f4cef41e7ba99b62edab616119dbbcbea;
defparam bigblock13.INIT_00 = 256'h597f0d98e8648ded608c2cbc6f26cd093a0c15027b771fa33e98c92b4fdb0367;
defparam bigblock13.INIT_01 = 256'ha8e87d1c6fc93a72b662a3471d83eec5dad28e360000801089cc1bf4dd65cb31;
defparam bigblock13.INIT_02 = 256'hb2b836bd62b938d934f60fd4200d5889000104005315689335bdfc52685d1d6d;
defparam bigblock13.INIT_03 = 256'hd65ebbae6696f417060e4ba89e7aa05dfd6b467bf4ed91c42fccbcb3d2abc89e;
defparam bigblock13.INIT_04 = 256'h2c10c2ce25efed17cdead72ce38657573377cd530f3c5c885608375bda1b8acc;
defparam bigblock13.INIT_05 = 256'ha25609162ea6e2a6e97e530d4fbf653ce6b5a6b3f30d051852e5ad95e6f952c4;
defparam bigblock13.INIT_06 = 256'h0580e6c01ea022342555d4f2135affff807ff800e32a558f922858cb7f7e8c83;
defparam bigblock13.INIT_07 = 256'hef4ac79e634acf1e27bb6db16f73854f402f27e24e66acd6cc0d400000538490;
defparam bigblock13.INIT_08 = 256'hac8c8a962b88df3239604ae6e41cd8a2dbe7980abf4af066290e99585a85d18b;
defparam bigblock13.INIT_09 = 256'h31ec49db0371ff807074fffbdee50a37aae33dac96d476d1ecb58368d8204743;
defparam bigblock13.INIT_0A = 256'h9f0ad7d4cd3ba3d89c38a8148b6d0087187e6ce635092e0c0d237b6723633bf8;
defparam bigblock13.INIT_0B = 256'h229938f9c0f53a077d1922a9d4e2a4c969533d027171b62cb7bb946d2896cd70;
defparam bigblock13.INIT_0C = 256'h0cc16f19aee68ca7e3a84da9aa0bab98db0074b62f659a601f992a147eb36c88;
defparam bigblock13.INIT_0D = 256'h83eb9541e5f388f8730e5ef590d2936e6c943b2134236f9e31fd6e6c91d1f0fb;
defparam bigblock13.INIT_0E = 256'h9025a526734e2c18641874cdce67b93d732f486d501627387b9450765824d4e6;
defparam bigblock13.INIT_0F = 256'he0ba4dc9fff9a2e6b70ef143a6ec69ccc91b833505c65440fab9fa30ee30a193;
defparam bigblock13.INIT_10 = 256'hc560680f428d092756884c32161a13691c91ef69a857fd0dd23be73cdf7de8b1;
defparam bigblock13.INIT_11 = 256'hfafd6c08393e95d2db2f9d8f2019f59f5fbee5af756d44b0d590d1839aa1a109;
defparam bigblock13.INIT_12 = 256'heb49b410292048177c9896aac967a7b7a8ef771fa796bdb8f2586e5d5b5f2b36;
defparam bigblock13.INIT_13 = 256'h9900a0fb7a10ec34dcd11551800474fffb7230ff2902c5da8e4d61474d9dbca9;
defparam bigblock13.INIT_14 = 256'h0011efa8ffbc1568ee3781614acc095850a36e5c9d12b728458c25734c11c608;
defparam bigblock13.INIT_15 = 256'h6c4adaaeb31c1c69eca392ea36efb425766e9df750c60c33aec3b4dfe391504a;
defparam bigblock13.INIT_16 = 256'he660675976791173d57448060149244063bd1800cde21f7028641a9d7c32900a;
defparam bigblock13.INIT_17 = 256'he337b9bd17efee58d5407bbc682f3b9d0ed36b029d8e403e292a16c9e5244d1d;
defparam bigblock13.INIT_18 = 256'hd497af967b9f0e0da351d4e8b6e1ac167581b35f231dac2e2745a6fd7d7d1d87;
defparam bigblock13.INIT_19 = 256'h3efb39b10c339c52f73debfad8a48c01798ef80807128b3002cb8c646d6bf2b6;
defparam bigblock13.INIT_1A = 256'h030e62b048009e9ba2360e7ea39952c43b68792a760ee120595fb994deb8fa9d;
defparam bigblock13.INIT_1B = 256'h08db42e6648639a9240b546c4bccd61795d7d74a6c9439c55d2232f2538a6134;
defparam bigblock13.INIT_1C = 256'h3e6bc42466d23f5d31f0ca08c55916a2ee3901158e03efbbe273a5d67627e5ab;
defparam bigblock13.INIT_1D = 256'h0d794c512804cd00049b682ee81bde690241000374fdfb7293ffc59bbfd9a789;
defparam bigblock13.INIT_1E = 256'h34ff00215ff4e9fb36739a7d167a7835681a57ef51ea548eef34bd1375608618;
defparam bigblock13.INIT_1F = 256'hc72d8b6a89b78f89ec9af1a9d5a1f8f2e15b968cb2ce45c70f71410cb3a2fffb;
defparam bigblock13.INIT_20 = 256'h494c7824b4f6faf5c97c62294a1f5df9ec14ded5969bb170200e046892dd036f;
defparam bigblock13.INIT_21 = 256'h166c582bddc25bcccc4a8907ddd2719378afec447f8f31134f7fdfa03033ac5d;
defparam bigblock13.INIT_22 = 256'he130bd0f87ca7508100336ebb79461dda0caf43d92ea54c2746a7d48d0974671;
defparam bigblock13.INIT_23 = 256'h2ce85ff97013bf88e2fd2c8746af41e93aaff63a321ffc18eed22c2a6478850d;
defparam bigblock13.INIT_24 = 256'h739542370321089a1a7a538c1828a92801021b8dbf5e25fb79e21fa554e7a8ec;
defparam bigblock13.INIT_25 = 256'h06d8dc28aa7b9c7111a248c34b3ef8601b57d95ba507c6cac5cb7db0490aaf22;
defparam bigblock13.INIT_26 = 256'h9a5f2330dbe01ba09f2a3d0f6e72880d7743d4ee3454b3ab0eeb0c87fed5a9e8;
defparam bigblock13.INIT_27 = 256'h9f92122044bd05734c4123a6992c649bc825861d5cd11e49000374f8fb72bfff;
defparam bigblock13.INIT_28 = 256'h794707af45ac0d2d2afa70f79d0e6d5914db24260000f765d40e09ff24166e64;
defparam bigblock13.INIT_29 = 256'hd78f20e684e0010027033f792809edf43cbe8beca9c972d894325d6bed9a0849;
defparam bigblock13.INIT_2A = 256'h78e508ce5ce22ee644ee1350bd6bd55afde46e8e012f45c30e52d5ab9fae170f;
defparam bigblock13.INIT_2B = 256'hdcdff9a447dfea609e931d54123a5028e18ec7b9d5b103fa55ca6d797cee2a61;
defparam bigblock13.INIT_2C = 256'hc8806732783ea5755edbc6db91241fd0a7398f26e1fdfff1bfd3b7f2b92f467e;
defparam bigblock13.INIT_2D = 256'h30600165cb163fd4276ed1c271a39bbb182e6ecda8981ac498544ac21ec8bd75;
defparam bigblock13.INIT_2E = 256'h9af8d0b255a983baa8f4e485b596cbe7960c8c64692a96dc18b1816f12905a50;
defparam bigblock13.INIT_2F = 256'h71b3b250b231c6b71e01ee44019d56f974e1cbe8d659aac22d50a1bbc1c6c5ae;
defparam bigblock13.INIT_30 = 256'h74f9fb705fff0c855f3920657ff449ddef738edf34811a96f6ddf46adce095af;
defparam bigblock13.INIT_31 = 256'h71d2141c6da8b3124b40433de96d0b08055c6619449b18258f445b3126418003;
defparam bigblock13.INIT_32 = 256'h9fdff73ba0e6c7fc8645aa5d59abb0513fab71b41ccc6b1e88db2700ef2e4da9;
defparam bigblock13.INIT_33 = 256'h6520659d94484280e916b142248c3693000a009006cbaad98b12ffe841fd23d4;
defparam bigblock13.INIT_34 = 256'h91947650d0ce3238a6747ccf92929ca4ebcd019cc40ec39895195e4ea736678b;
defparam bigblock13.INIT_35 = 256'hfffffdbf1dbfbffdfc865fcd14d2b7f383576e60de716223703a4d74c716607e;
defparam bigblock13.INIT_36 = 256'h46510010df04b875f4a6824ce10f1a3044bc956b0e3616d20000facaa97ffa9c;
defparam bigblock13.INIT_37 = 256'h1303436104561b8e20000120daca0202fe3e4de41b4037be43855c06045fbf04;
defparam bigblock13.INIT_38 = 256'h2a3ecc4cdc971b55ccab4ea1068ffdd40411de498d2d90c35d136996a864b96c;
defparam bigblock13.INIT_39 = 256'ha47b6f7f8991fe4d61f7faa0a9127edeac73f970dd7b6d6aa06bea69bf3de7ff;
defparam bigblock13.INIT_3A = 256'hd1eb41da02d2fc807274fffb36bd2b8d00294640e200e7f99732fd1f3f96ffe5;
defparam bigblock13.INIT_3B = 256'h0c4509e52c947c09adf04c6213ed609ca5546ac7f1257c4b24ad9b5730443d40;
defparam bigblock13.INIT_3C = 256'h0faf66ecfd871cf94083ba0340a865438161ab6e5465e428cd39bcf4ce9a7f45;
defparam bigblock13.INIT_3D = 256'h9e4cd9ca914b190f2d15e2f34ee2a3650947300217065ccdc9ac8aae9faf7c92;
defparam bigblock13.INIT_3E = 256'haf4f19cddd8fbc0ac4267273b5357fe6422d8dc08cff1c01a432e717d714c1d3;
defparam bigblock13.INIT_3F = 256'he77fffd1fd5b86ffbffeab1adfbf14743fd5f38f03f34d0b38a34be9781e9efe;
defparam bigblock14.INIT_00 = 256'hf0a230e09753876637605281ded6cc93e35d7256a0333e301568fceb8e76ee5a;
defparam bigblock14.INIT_01 = 256'h364a280096ad4000e65108c13e1051fe8a37e800b870678f1330b50560262a5c;
defparam bigblock14.INIT_02 = 256'h80ae8b150ade681f075470e49e88bc29449fd897a78622724a7387b6bcc31d59;
defparam bigblock14.INIT_03 = 256'hcddeb1e4a7d09be64ae00d684f1e0dbdd21a85e09d158fa911b172a3d7f9248d;
defparam bigblock14.INIT_04 = 256'hbb6a2e0454a0692f5f5b02d1ff007274fffbf63ac6fffffc51d99fe9a9ea9ee7;
defparam bigblock14.INIT_05 = 256'h36d480607a205815e1474269cdff3ed0b4b492ed40ee2cfa6da6e907c20a204a;
defparam bigblock14.INIT_06 = 256'h7430ef9c5895a02ac6c0135599f710673eb55e1aad0d5b0b9855933dcac16e35;
defparam bigblock14.INIT_07 = 256'h0fdd8bd915c2cb0f070f5586e660623a0a0d000022e0da01250de07433fc1bf6;
defparam bigblock14.INIT_08 = 256'h99fb750d393554b0dee8fcfb877e173022376bf6be84057bae8386bcfdeea45c;
defparam bigblock14.INIT_09 = 256'hff855367576a955f322916cd84ce67eb1e7ad105650748793485b88863a77b01;
defparam bigblock14.INIT_0A = 256'h68fc6d12dc74dd3b6db5349c00075be09945be99d5fe9bfa41ddff90e3fe9fff;
defparam bigblock14.INIT_0B = 256'hcd68502ab32600100502500150107c80797745df96b646102f1bb7a458dd02ae;
defparam bigblock14.INIT_0C = 256'hbbaa01dc0823bc3eeed988b29f4fe05aa449d498fa2adadf1975a439c76f6a45;
defparam bigblock14.INIT_0D = 256'hfeef3c5491be3d110694cf28c543d32d3596781ac424abff9bd2495be7d1cf72;
defparam bigblock14.INIT_0E = 256'he55b6e4b18ab9b8a2f643b7269895e5c02effc807274fffb8e90bebf8269754e;
defparam bigblock14.INIT_0F = 256'h6a2038db892d5562c9151010ffe6fe8d20bfffa73708288192ee60bab1527144;
defparam bigblock14.INIT_10 = 256'h866c1048800219173b1caabf471f6c2294de0e76353148976670d764e56abce0;
defparam bigblock14.INIT_11 = 256'h70f1fd9b0264c6e60ea2c1f46e1fd569f098eaf8f354e4338e313a7a402edc72;
defparam bigblock14.INIT_12 = 256'h3840a5246c8297efd7fa6a25fae0df3370c3529a074e5c09bb95997b156b1f86;
defparam bigblock14.INIT_13 = 256'hf77770f0e887f735814773aa32ff100c4d6528e61e7a180ae050b596d68b9c6a;
defparam bigblock14.INIT_14 = 256'h189b1dcd9b6fd62bc8b204adb6940371fffefffffffffffffd3ff9f709181a16;
defparam bigblock14.INIT_15 = 256'h4f93a995a8546d32002210004da6f9a4abff7ace31c94d00dda5f6930f7ca368;
defparam bigblock14.INIT_16 = 256'h8d356840d946864cb501f51b71bb6349e5d6263cd66945961706233b85c60c4a;
defparam bigblock14.INIT_17 = 256'h7a7f30be738d0e6b6b631e0b250ad0cb119fa83a5abfbed21d3ba904e990172e;
defparam bigblock14.INIT_18 = 256'ha07cacf16ce74d5b900c1988db6a23422dd8398b5fdb033bfa007074fffbcfb7;
defparam bigblock14.INIT_19 = 256'h720402da895130beaa550756ffea1c2f8f1cb072f4fe3fa7fda5adc98c910aed;
defparam bigblock14.INIT_1A = 256'h1448765daf6ca9060fe321710400370bab2907a337fa07eab61ebfad695c1500;
defparam bigblock14.INIT_1B = 256'hfd5352812455cc10dc356833ec98d08fb45411839c96aab9c2b440702c75d3ba;
defparam bigblock14.INIT_1C = 256'hf3145dd2d257ce8820f4fa8e83ac15de80b1f456b3b7e9cc03a7203f3410bca6;
defparam bigblock14.INIT_1D = 256'h9c8d0080fffcfffffffffb45f395e9bbd47f9fffdda4d9ffa55ce8750f520772;
defparam bigblock14.INIT_1E = 256'hf7aef33e77f08be4c60bd9d97514559ea984ca981928868d46cb705cbcbea550;
defparam bigblock14.INIT_1F = 256'hc50b67ac88fb3fb4ddaf1bd1f9fefd651d7333d1f37c73c5968e064f800074ca;
defparam bigblock14.INIT_20 = 256'h883652c16b6797db5deac0856c94dd0cdeec306ba54ae363295b6cd72df911e6;
defparam bigblock14.INIT_21 = 256'h74fefb729fffe5ffe7fffff1b06363a896ea92ece50caf3b1d59b92055ec32b6;
defparam bigblock14.INIT_22 = 256'h9157c32decc8840a54c067ad07660b25e942332502db88248d2f5989af498003;
defparam bigblock14.INIT_23 = 256'hb45ac4b6b3c69ddf0693dcf20d8c844aaea2216cd7156e382a02a7d02cada819;
defparam bigblock14.INIT_24 = 256'hd501b37f415c48fe65f276b312d800cc010000024610179c0485ef6a194eb644;
defparam bigblock14.INIT_25 = 256'hebfa39ea96bc52d4aae587af1937de48b24209165bc2cd2bc5e8aae22505a186;
defparam bigblock14.INIT_26 = 256'he64f10d34387d356764c0f4d5e5d2b21edbb5d1de928791e6989d2d79a0d37ac;
defparam bigblock14.INIT_27 = 256'h40b9ce205101c6db400dffc0ffffffff68ffd55d926afd9f7d4fd87765ff5082;
defparam bigblock14.INIT_28 = 256'h01348000265c6e75f96dd7af01f25025bf38bc8f30256d631725f63e9793461f;
defparam bigblock14.INIT_29 = 256'h7d672d01f672242665cb53a7a78d4f4a1338c44f5434b56832980223b92715c3;
defparam bigblock14.INIT_2A = 256'h648a5daa6a1ca40235a25a7a8bdec886e9a0200779cf3d3a89cc6e22d4ec4220;
defparam bigblock14.INIT_2B = 256'h58914e49800374fffb727ffff975757fea327a3d455bae6253eb0cbbba172ba8;
defparam bigblock14.INIT_2C = 256'hf8d3f3d677ff60ffc7956c4c948b514047b125620c11e9501731a2db5026eb6c;
defparam bigblock14.INIT_2D = 256'h3fb0767cad106a4a564f6a50d816951748dc233c244eb1750815db4b01b8ff8f;
defparam bigblock14.INIT_2E = 256'hcd3276c068d5265f6b0cfbac8b315713b97e0edb1e650007010402f6d43da5c5;
defparam bigblock14.INIT_2F = 256'h09d56b97cebc5cca14753910b082f6568fabf614fff44a9845c6d905b9a99e74;
defparam bigblock14.INIT_30 = 256'hf8f177ffaed4c7bfe8c44f57b9c4808b230ad4933d8a817aae079d93bf034cd0;
defparam bigblock14.INIT_31 = 256'hbef98d50b8dbffe0ffffffffffffffffffffffffffff88fff437f943f2f69fa7;
defparam bigblock14.INIT_32 = 256'h0099b1006232db5cf0af19e2fc58ee9c2cadc9e3e2920b355d89d5872829cb39;
defparam bigblock14.INIT_33 = 256'h59bc35a96272d20a85dbc6cfa957262104572bb44e0dee4baf215b4c29f6af52;
defparam bigblock14.INIT_34 = 256'hec59c0349cd95eab0c8bfd2887dfbe7842262284ff40775321688845bfaa60ec;
defparam bigblock14.INIT_35 = 256'h62dba027ed1658c94a41800374fffb72ffff336f5ffe480eade54bf9bc7a1e77;
defparam bigblock14.INIT_36 = 256'h512a0724f52cdfabf52ce7ff084297a26c4c900bb4c047ad3f620c2deb381725;
defparam bigblock14.INIT_37 = 256'h0c00088267f6c762927ca38269bce9fd4a32c8ca5837bd4f708ceda3a2e3ae8d;
defparam bigblock14.INIT_38 = 256'h381dc7d028cdbc6780a41f55f2e1a2186f5da8d1934bcf68e84d399001640021;
defparam bigblock14.INIT_39 = 256'h9b26b031411f51d2caa713421715fcb32e5d5b62f085771c16d5f28bf4caea48;
defparam bigblock14.INIT_3A = 256'hc8a23ffb157f1d9b7b94f0d55ef11a11ad77b410c4a06a70a10aa9468ed5ae57;
defparam bigblock14.INIT_3B = 256'h025003c8162d048426960b72fffeffffffff4fff1bde6f35847db668b2e79953;
defparam bigblock14.INIT_3C = 256'h4c210c0b0d4c0110004150518aa00bf9e8bb161cb480b721cdf4ad4cb83186b0;
defparam bigblock14.INIT_3D = 256'h908eef25888d8506dbff80108624f7ac12e17d6042d21f557fef465a795cab64;
defparam bigblock14.INIT_3E = 256'hf8488ee3b221302437b4bda3cfada1e41b8dfd9c7eea071fe9274c04bdde7c45;
defparam bigblock14.INIT_3F = 256'h0b69aba0133022db30230c3dd8b39b41800374fffb70f9ff4d7f5fd06cffdffd;
defparam bigblock15.INIT_00 = 256'h93a46b0fcae302212c889f12db6cbfecfe9d087fc7966c4c8d0b54c0a7a53f62;
defparam bigblock15.INIT_01 = 256'h00120040000028021d3277fc3d22cb7e9a0544744c1c15de56ca185ac48581b4;
defparam bigblock15.INIT_02 = 256'h524512b9931f23c1db736623de33b13156ac161ca4874fce263d904676b366ea;
defparam bigblock15.INIT_03 = 256'h24b2dd4806265426fd4ac7b53d3b87fef6b77bb5bb8658f1cd500622d6a97aff;
defparam bigblock15.INIT_04 = 256'h153beff4ba9da2611afe576a1413daafcff5f409aa7040b91b9c21e8d1a8a772;
defparam bigblock15.INIT_05 = 256'h3eab43544c8d824360c2eb82963971b6001380002008da0674e5bf20e3c17ff1;
defparam bigblock15.INIT_06 = 256'h8c8387f284f4028a2000020122001a20acb1fe667b4e6ebed1bb79396f419513;
defparam bigblock15.INIT_07 = 256'h2360e9d5a4c250e07dea6168abc859d493ed8fda2f3474f9ae1191b2f341ae0e;
defparam bigblock15.INIT_08 = 256'hb2147bffffbc3dd8503f32a0278f1d7dc048513e2f2e0e1b8226a11d195c44ad;
defparam bigblock15.INIT_09 = 256'h48852c5566e6b9754a0b1927db33220246a8c1ed425903a7ff807274fffbfffa;
defparam bigblock15.INIT_0A = 256'h3767e51a240064b18d6226e300086068e65829aca5bfa90f17fcad90dc918b6c;
defparam bigblock15.INIT_0B = 256'h859120361161200800000140129b97fc5268b51b80b3770745cfc2a3e523595d;
defparam bigblock15.INIT_0C = 256'h348c9028e738c1aa1e8810ba94232d4ec9426603ed296d71304406d90c04a21b;
defparam bigblock15.INIT_0D = 256'hfe8c1afefacc56319ed6090065697776f93bf2a0464bbc78806b12506bcfe3e8;
defparam bigblock15.INIT_0E = 256'h7d03e8a5dccb5126767d2736851bd6966b1ab91bff01fe8fafeae9fcd0bf7fff;
defparam bigblock15.INIT_0F = 256'h4f60c1e126ee5cee52d1cb5a1646d6579083098fa1920400c1c2bd9c7e8520ed;
defparam bigblock15.INIT_10 = 256'h3abd47996ecd80372885ec72a51dc7e762e4bf1a4fb883fc06cbfd3e43baec66;
defparam bigblock15.INIT_11 = 256'hb6e7a16a91d03d278a37465ec9655aaa7a19789c4354c53c4bfac8adc9048589;
defparam bigblock15.INIT_12 = 256'h7274fffb51bc5fcca7c5b15bd937d94f389f3d03ec99262991f3dd5fda26ef90;
defparam bigblock15.INIT_13 = 256'h2d51e8938aec408dacf467a76505200b2569db3d26c23f18e1ed4f59038eff80;
defparam bigblock15.INIT_14 = 256'h9bb442df3ae8c4fec711d41a5e6130ebb06da5119c6d0104608437dd14ea1a0d;
defparam bigblock15.INIT_15 = 256'h37b1240b186ff69b14146296990e4001006bda002a9408caa9b42756fe69e885;
defparam bigblock15.INIT_16 = 256'hfa782d67077e1b6bb6aeb74b0bb6824c7cd8161511e4ef5b52c5cf92155c662c;
defparam bigblock15.INIT_17 = 256'h26a01b2609ad93ddc4519b62fe36bde52635e4c2aea5d5c7888bae316a60bb6d;
defparam bigblock15.INIT_18 = 256'h0044bfe8db524f754e830281db852c191fee817d79414ffbe81ef7d57de97d77;
defparam bigblock15.INIT_19 = 256'h2810a6608dbcad8f0392e236a64afd60aa83660124963673d4a113216db510e4;
defparam bigblock15.INIT_1A = 256'h8446262396c14e780e01d8e903f70bd49b2ba51589a182c742dc70ca44860000;
defparam bigblock15.INIT_1B = 256'h4d155ae33dbc51b98a209af82108d0045c3ad365defe66c8cc7698e010fae58a;
defparam bigblock15.INIT_1C = 256'h415a02b8ff007274fffb7bdf5119b7b875498224ab9f46f8ec7c090ff7df5545;
defparam bigblock15.INIT_1D = 256'hadeafd20c6f7a4481c910b6de095317368a6893d620f24c7db431c825480612f;
defparam bigblock15.INIT_1E = 256'h08c499a89c5ba5de66525a61717c942db6fba1056d60b8dc0168f24aa63d889a;
defparam bigblock15.INIT_1F = 256'h5487fe4053280e1749e347bfe55e98d95b59be3b00060042829065e0f5aa2db1;
defparam bigblock15.INIT_20 = 256'h4fde7acd2aab1ec14ddabaeb6c98c7bde28b2641bfb2341fe339722fb24add69;
defparam bigblock15.INIT_21 = 256'hc673346edddf1f12937bb30abf69363327b9149abc2ada50a30716755642f968;
defparam bigblock15.INIT_22 = 256'hffffffffffffffffbfff70a15653d402e24bfad22f0cbf8fafe6246b65f5ed9e;
defparam bigblock15.INIT_23 = 256'haf7d8044b9d2128c6ae7da8211b4b5b38e8c0c0cc8323a596d50b7240140ffff;
defparam bigblock15.INIT_24 = 256'h7529e6db21319bb56b87dd1afaa523a573e9a8a60c2501590000b134e718037e;
defparam bigblock15.INIT_25 = 256'he528c1175a038f272196a039155144106cfdc48a8407274e4e7085bceb1bb650;
defparam bigblock15.INIT_26 = 256'h20021798c9eb485a0383ff807074fffba16f77ff7e554efda163557f43935385;
defparam bigblock15.INIT_27 = 256'h225b4d0083879a9fbfd2ca7e89695cc50aede088ac536ae4953d644c24c7ab5a;
defparam bigblock15.INIT_28 = 256'h63851da06c803f8a93aa62ce4bd7188c58f5eb48547a95eaf28fbb78aa1791b6;
defparam bigblock15.INIT_29 = 256'h417e801054dda0df5f96c28726bc442f91012b236a5796078aab001009800000;
defparam bigblock15.INIT_2A = 256'hea464d518edd07c37df5b94e9b6331013c3f42eb06239f426a385f51623b9ade;
defparam bigblock15.INIT_2B = 256'hfffffffffffffffffffffffffffffeaf4ff4f6fef5375229ddd93f92f7744224;
defparam bigblock15.INIT_2C = 256'haa96161360ea0183ec39b4b0402a4264b60f8f1199c883eab582dc6d0124fffc;
defparam bigblock15.INIT_2D = 256'h5ed166fcda7301fdc955589d34a60abdc9be9a41257b176e5080e4a696eef292;
defparam bigblock15.INIT_2E = 256'h567fa4c74f46060e5d9ff3511e5e1ef7fee204189db540eabdd95840d6289bca;
defparam bigblock15.INIT_2F = 256'h14c3a86cd256e664fb6ad4c86de03e9c79db129c542abd689ca15fe9e0f5d404;
defparam bigblock15.INIT_30 = 256'h0a752d1e373182dbf823ec5a59b1d048800374fefb72d1ff13999c1b3ab3f655;
defparam bigblock15.INIT_31 = 256'ha13d36da006ed00159cfe9fff2a0a67fe4a498afc4896cdc8b8bf64067a00566;
defparam bigblock15.INIT_32 = 256'h9590836dc0114ac65ddd7e508c6e60c079c23ac2d52190aa38a5cab4f4bec81e;
defparam bigblock15.INIT_33 = 256'h95ca193365b6fcc3c913979a1fcdd05ea9118863a0add473448d49aa54e5bfb4;
defparam bigblock15.INIT_34 = 256'h9f2aeb18afcc0fe97beacca9eaa823668e604f99c6f8d4f213871ad315e506ff;
defparam bigblock15.INIT_35 = 256'hfffffffffffffaff57d77f93f949abef8a40edfe17ce37adac2373be8dd71500;
defparam bigblock15.INIT_36 = 256'h568f20a4d10c06ad181b8d225925d212a5511c6dff81ffffffffffffffffffff;
defparam bigblock15.INIT_37 = 256'hb8ea3e50c52e1ca43f49c67a025c5d0f190af1102c4212de69d3ed04d97fd726;
defparam bigblock15.INIT_38 = 256'h565f63154191619187d2d7bbb60cb9bf1166f01a8a562533894121444b36b236;
defparam bigblock15.INIT_39 = 256'h6fd5532b79bb273e4c9b52018a6f7d6e254b30d982d94d56d94e9032d3600e59;
defparam bigblock15.INIT_3A = 256'h55a027ad3d660dbd2b80372442db30258b6dd9c90e32800374fffb7275ffe91c;
defparam bigblock15.INIT_3B = 256'hee013103220a1a484a0806c3b6d6037157d2abedd9f6ff2889dfc31decdc848a;
defparam bigblock15.INIT_3C = 256'h84999cf8a8e3327f00110400060ada22e974dde886a1c5e14eefe423b6b60135;
defparam bigblock15.INIT_3D = 256'h9a11ddc962dbafb08b7cf52f780835be87efd30b7456fdc1a1d4699e90ec2da7;
defparam bigblock15.INIT_3E = 256'h77fff5775dfb7634bbb7d475d28054bcbfa64074bfe0f9c4c100a00115aa205d;
defparam bigblock15.INIT_3F = 256'h0803d31a69f229137fd0fe00ffffffffffff5fff7dce0f3557fa5bbdff92f96f;
defparam bigblock16.INIT_00 = 256'h10cf755148658694117ef1c1f1d025a5fbf80b8ee41a53e438223ca3600b9383;
defparam bigblock16.INIT_01 = 256'h6bb4ac914bce1589eb2452f9c3e96817b31e2b87796b32ca000096400be5c463;
defparam bigblock16.INIT_02 = 256'h3f7e2e20efd9a80d488cf67646f000d56b2cfc864da97634b45b2ef85d8477d7;
defparam bigblock16.INIT_03 = 256'hfb72f5ff6b7ffff58a96fffdff98696f8dda793201f5c8c4cae52fec3c4a9340;
defparam bigblock16.INIT_04 = 256'h94946c4c908bad0007b107624b7de8901331e2bb9024ed56d8898948800374ff;
defparam bigblock16.INIT_05 = 256'hf3969be5b3068435b9adc6310b8da8cb02bcb8d4028de64aefe32979fd91f8ff;
defparam bigblock16.INIT_06 = 256'h4abc2f72051b918ddd190dad818d04d482006a204d1eda666a5d3fbe10ad958e;
defparam bigblock16.INIT_07 = 256'h5893b9341c2c8ae80f847520f2f01a1e57318b5a7625bdc9a9e31111ab859976;
defparam bigblock16.INIT_08 = 256'hc015e930a467fa680ec617903129feebfe9089c110aaa9dd8506371d23761227;
defparam bigblock16.INIT_09 = 256'he040ffffffff970ededf60694c207f4d60c2fa7e0ab3d7e8239bac2327ad674d;
defparam bigblock16.INIT_0A = 256'heae142dfcdf9187cc1786a5a781e264b0ceebf503253c5c12bb50a7a8da986e4;
defparam bigblock16.INIT_0B = 256'h25dade95b48dff46aa43555b26a0040bf06bb948333f585300000012c0006800;
defparam bigblock16.INIT_0C = 256'h88d2fac2a6128769a330c5e350dd423ed8c886229bb21c2b6125658e9a0e58fc;
defparam bigblock16.INIT_0D = 256'h0748800374fffb700fff4aeebfc5fff24656effffb20be6b2a1f1a54a9a6fe63;
defparam bigblock16.INIT_0E = 256'h2afd320ea8ac66346c8c8c8bf84867a477640c216768222504bb1030e23e5919;
defparam bigblock16.INIT_0F = 256'h17a74a34066bfb416a347c1977ec25af17ad0bb89141db6b0938c0000ac07dd1;
defparam bigblock16.INIT_10 = 256'hd6f1636515662d9410eec2e991c0986b6eabdc61400101009047f68cd776a7e6;
defparam bigblock16.INIT_11 = 256'h1ea6870af3f3c630da25ddd9a8a422913c3bfbb065be9e52dd7a5c33bb5a0b54;
defparam bigblock16.INIT_12 = 256'h3eafeff7c4ffeafc3357eaf7f65d09e6f40c694f17458625bab82b286af30fe5;
defparam bigblock16.INIT_13 = 256'h582c50dfcc5e541b4af99d17620c4094aa7a71c6045bbfa8c3a25bba15ea2852;
defparam bigblock16.INIT_14 = 256'h2dd1d68b76614db4a54209b6ca6257d2d33c01510010e4000794b3e75ab002d7;
defparam bigblock16.INIT_15 = 256'h605574172e129563f8ec0490ffb53d856844c0b12b6080105b03a5774fdc6ad8;
defparam bigblock16.INIT_16 = 256'h113db0e130507c4e8a2ca89604812a85240cbda206ac700a496f9486962322e7;
defparam bigblock16.INIT_17 = 256'h22a23d58b1ed4fd9038bff807274fffb3a0b401470f04aa13c8134f512950c7e;
defparam bigblock16.INIT_18 = 256'hf1f77bf547eadee11e2a173d2da0e8c40b6c008f3d5267a6c9050e0b1928db37;
defparam bigblock16.INIT_19 = 256'hd1304ae1d8d12541072859cc1b6d51b90007d7001bb6633d64b9f14f69cdbdc5;
defparam bigblock16.INIT_1A = 256'h90e5b468bf6d5a726247e79ecb8719162babaa5e615c32962461000e01406ac3;
defparam bigblock16.INIT_1B = 256'hdad37144acf559660f5b6369d7ca0f5a2dd46914d6ad218be5da66b3d05910a8;
defparam bigblock16.INIT_1C = 256'h331194cf555433b143c31ec0aab44bb90b3ba0c36d010a5cf65cb366bca55743;
defparam bigblock16.INIT_1D = 256'hc080ffffffffcbafc495fc64b8ff455df5aa558f67f76be91baf319ad6b03d6c;
defparam bigblock16.INIT_1E = 256'h47db7da528fe01c82040000235b25ad91fb8b7c620384513882a6a88c91b0371;
defparam bigblock16.INIT_1F = 256'hf5f559284923d3b449bcb9d9b9f7b881dcfaaf6f2cf724069102d201ae633623;
defparam bigblock16.INIT_20 = 256'hd913851d75c2ce973553d2c77f0247d39afa2431f0c0aa3f55f6784b115a35eb;
defparam bigblock16.INIT_21 = 256'h66102507db571ee26d28c9e9485a0311ff807274fffb4398fca2277ab9d5ccf3;
defparam bigblock16.INIT_22 = 256'h896e102092c727d6fe9122efa7f4ea3bcdef0c89683305adc853b1096b47295b;
defparam bigblock16.INIT_23 = 256'h040b0022cf00054447fd67e520446da9c8d6387ec8363d735c441ad8566646da;
defparam bigblock16.INIT_24 = 256'h2b656b313923eca49e6b666c8d458d8a6bc8ab8b1f38ae3bd4f82379e366d533;
defparam bigblock16.INIT_25 = 256'h4cd61d1f01a1cccbfdbff532f9f1de8b9e2f19f31eabfc1fd2fdf2beaef52178;
defparam bigblock16.INIT_26 = 256'h8148bd0417b95d2e44b75b6f5e3e9422a0b832f79bd356570c37a054bbbd8fd4;
defparam bigblock16.INIT_27 = 256'h97d936b51b8efff0ffffffffffffffff751fa6347523916a5be1812d4ffa58f9;
defparam bigblock16.INIT_28 = 256'h32cc10000c95990bd07b67484c9eaec81afdd8fab0ffd68f5dfa060c25a838a4;
defparam bigblock16.INIT_29 = 256'he8af5f2422679426ac36a1529a3e63ab7f1c8216a9e7c96243138fe5b51985b1;
defparam bigblock16.INIT_2A = 256'h7e99d555784084afb229913d3c2681ff54f1058b4415c733d53164c9625004fe;
defparam bigblock16.INIT_2B = 256'hacb56b279d5b044c0cc64b5a15c14628b1ec565a03e2ff007274fffbb5baa43f;
defparam bigblock16.INIT_2C = 256'h0e18641513e0e0c7da446e36c5404fffca7fdbffff43226b1ce85c838b6d6078;
defparam bigblock16.INIT_2D = 256'he954c45b31b006b0480064008502391f3f5c038d4768fe0c9aaaa19717ae3751;
defparam bigblock16.INIT_2E = 256'hd0665676a18030ea719d286406a4eead766850dbad29302ce880f4d33c8f20d2;
defparam bigblock16.INIT_2F = 256'hde25ad5f04930d8cec846e6130beae83f1d77ea318fe01599878c603bac91d30;
defparam bigblock16.INIT_30 = 256'hfff0ffffffffffffffffffffffff27fffc89a6fffffefffefffdfe3e917f7ebf;
defparam bigblock16.INIT_31 = 256'hf9fd8eb99578abab752327d17f626d238759e45a4311406a4ddbd30a8e460403;
defparam bigblock16.INIT_32 = 256'h376a3c37e9a5503b8d64411b49d32f199f8e18f3a60bc000202582753d7a1105;
defparam bigblock16.INIT_33 = 256'h2f3983e589253e3cce15217990e9fb479b5cc182726215180cd4ec64c7b196da;
defparam bigblock16.INIT_34 = 256'hfffbf975fdff37a8df537313bd73f39487a43d9bb736dc8a9a58a1fc4eba8b0e;
defparam bigblock16.INIT_35 = 256'h8c650b6c4087b14d64476923900a31e7db232282471811ec48d903f4ff807274;
defparam bigblock16.INIT_36 = 256'h6b55a539d8a1ac40b6fc839b54c838479458db502e38acb8f9efff397f5b9cf8;
defparam bigblock16.INIT_37 = 256'hd33c1891ba413fec4f068cee4dab3aef100043ae7e755163667e184bc551ab2b;
defparam bigblock16.INIT_38 = 256'hffb29350062e4552ba8d895430a9bf4a23b591b3f2c40dbd51fc32eb8de3234a;
defparam bigblock16.INIT_39 = 256'hfd5b03359a84c39f325ce8202d518e84b6c702a1705946fd53c7133f84006032;
defparam bigblock16.INIT_3A = 256'hd2426e36ffc1ffffffffffffffffffff883f9577eefd5677fb7ee367fcef538e;
defparam bigblock16.INIT_3B = 256'h672078f90c94ed84a2a6b990add1d9b78ee98ceaf0eb496984d958f8e3b34885;
defparam bigblock16.INIT_3C = 256'h4d158e40c29357f00521088b60352f5382d8dee654d7c4a2775a7ba211c80000;
defparam bigblock16.INIT_3D = 256'h0a5a994373b2abb1d075b29811943a2563851b33e452690e3fbbc62006c99a7a;
defparam bigblock16.INIT_3E = 256'h0354ff807074fffbfacda5d7cc13b75a24bfe9296b3950b210252c89e9c4a5e5;
defparam bigblock16.INIT_3F = 256'h297f15bbae084cc78b6cc091adb462c7e905900b31ebdb1726e25482b1f85e58;
defparam bigblock17.INIT_00 = 256'h821dabb43b401e404d0bbb34946eb87c4fa28a37b4c1dc6d4800f133b2b3ddf5;
defparam bigblock17.INIT_01 = 256'hee0d2ace78c1a00b93ae8d281a7de72ba6b9c4ce000401401d127f349b5dddd4;
defparam bigblock17.INIT_02 = 256'h44ffa1342fd6b62932fd362d3fa2473d8f69970747ece88be9fc629db4c3a3fd;
defparam bigblock17.INIT_03 = 256'h6df96ead301b61f7236e199dfa4aecaab4176e66b22fa648a21e8930ce32935d;
defparam bigblock17.INIT_04 = 256'h609726a8abc45b7f57d647beddda07fdffe3ffffffffd227f46c2797feba6baf;
defparam bigblock17.INIT_05 = 256'h5120802087cad02675ffffb18925303807f21683d419d080f13fe7e7d6383153;
defparam bigblock17.INIT_06 = 256'h579a598ab45cbd48498e4df8a35e4937e224512f5caa26b929195f15d36d010c;
defparam bigblock17.INIT_07 = 256'h547245bf417e8e82074141f2f116cd3bc1b7c7a27443f97c85100524a426269d;
defparam bigblock17.INIT_08 = 256'h2023095558936a48800374fffb72b5ff91710d129c187f66ddfbf29f6ffffffd;
defparam bigblock17.INIT_09 = 256'h441b636c441d5ed845549018c2b56c4c838bacc06c3105620c85e7581325c2db;
defparam bigblock17.INIT_0A = 256'hc953f4111c2fecb798f1113c42f93231280817101f543062e6a9371c90424b33;
defparam bigblock17.INIT_0B = 256'h20033118d8d55a901086f11da3c0603be58453a40dd4960a42a0001100008f22;
defparam bigblock17.INIT_0C = 256'hed283be49217cf4878f826b638040688de3d4ce58812090bb4643f7a19a8c595;
defparam bigblock17.INIT_0D = 256'hffffffffffff8a7f83e0dbf839ff09fba7d195d3f6bf1a5b2faafacb2b064f28;
defparam bigblock17.INIT_0E = 256'h10eddab603f2315bcfabd3431d3ac9140ea91d1a2b2a6b14da626eb80000ffff;
defparam bigblock17.INIT_0F = 256'hdd0dce4e0902365d5e4b02364c51b0592081e0528af279e16829000608049472;
defparam bigblock17.INIT_10 = 256'h17ff4ad7f59b217f3446c373ab7bee24888c275ac35d4c63e2f9e98576d52070;
defparam bigblock17.INIT_11 = 256'h47203630463d59f5005cd289cdffe26cbdfc5b0819fd6f26c6d8ef76418ae964;
defparam bigblock17.INIT_12 = 256'h6868323cc49b582ce96bd9b13b4f800374fffb7270ff65ea675450b45e9963df;
defparam bigblock17.INIT_13 = 256'hb6ba1c919e826ce8c41e177aa0895953a1d1911decccc3934cc0e7b103660a21;
defparam bigblock17.INIT_14 = 256'h00260480a694e4e8c2c2bdb50720e21584158ed53d16f35651a622508d452369;
defparam bigblock17.INIT_15 = 256'hc6cfaee6692b11e15b621573d72292a4c3b34799783a4520326975cb00183400;
defparam bigblock17.INIT_16 = 256'hefb8de1d2a9efa443affbc3814a77bf8b62e1cff7efec5e5d8aeee19af5fd0f3;
defparam bigblock17.INIT_17 = 256'hef52d21fdeca826c84afa9f4732397b913b455be1144bfc9f4f7049276d41ee8;
defparam bigblock17.INIT_18 = 256'h83172f173083839c5548c6db520d0002fffeffffffffffff2fffc74a7328bf50;
defparam bigblock17.INIT_19 = 256'hbdd921483007e2cbf70d1ed1a52c12d4031d00000bb07f08fc9c18689341b916;
defparam bigblock17.INIT_1A = 256'hac1cab5584c71d1fbbedcdae856e561fe9bba9c55d72b3b50033291a77a2c5db;
defparam bigblock17.INIT_1B = 256'hf18435c05cc16c33688af9d4575e94d403055d4aeba35acf6f5b0396f6b5deb9;
defparam bigblock17.INIT_1C = 256'hc63d23640ead654a272542db2020e953d919ff41800274fffb72e6ffdecc71e6;
defparam bigblock17.INIT_1D = 256'h6dac16e4280026007a5e95b195fab9e48232fa75b10cc842919d6c8c820b53a0;
defparam bigblock17.INIT_1E = 256'h55a55816350c000280800910a7f2dbf4031ff906c7a47aeac1b00c9dce93daa8;
defparam bigblock17.INIT_1F = 256'hf678520b095d818f133ddef59ca113d9a69f37cacdd3fdc2bb6037409c57f2e4;
defparam bigblock17.INIT_20 = 256'h654ec0a9543499a9714872ae235ad5747fe514d41be3d9c152596fdbf34bad9a;
defparam bigblock17.INIT_21 = 256'hffff390fe2c24f44fc58e21711d99fbb96057e884cba9a3cdf7a476e8f85574b;
defparam bigblock17.INIT_22 = 256'h424274e0f8451a2f73aaa4b5b5996042091e0761f2e76244358cdc8e2102fffc;
defparam bigblock17.INIT_23 = 256'hdfc4d4ababf4bbb66e7a7b32a762ba28cdf844e4c8dbd482ca78011b800008a2;
defparam bigblock17.INIT_24 = 256'hedf101a4783447f587a49dbb5e34a0d47b73b7a66fe62e0b8d48195f99717c61;
defparam bigblock17.INIT_25 = 256'h1dfffd058593a884adabceeedc75d152c6ef3c049ff896b5cc8bc504ae58e5f4;
defparam bigblock17.INIT_26 = 256'h2de8700b5e60e620216e0d5d48387a0c41fbd81a2f445be99f41800374fffb70;
defparam bigblock17.INIT_27 = 256'h65c6ec588533d6abd97236d60b8e38200d003d70cde8aa7ffffde51d403f648d;
defparam bigblock17.INIT_28 = 256'hc4315acfca3331dc24b800c4000000002f4ae1035bb3fedd97a85412f1a8953e;
defparam bigblock17.INIT_29 = 256'hf08d83cc8986b80d54db409f97f0495f40a2935d3151924313b484aad85dc1b6;
defparam bigblock17.INIT_2A = 256'h808ef46589893fc7dceac048c7c03914ccf928723e2a667f7fccd84999d1ce60;
defparam bigblock17.INIT_2B = 256'h8cd5ad17d8eaeb54db540dc6c100ffffffffffff4bff961edc2d2dfee5fff137;
defparam bigblock17.INIT_2C = 256'h595ce86885589b2e135902480000f8b98c83ba70e81af941b32dc08f2706ba4c;
defparam bigblock17.INIT_2D = 256'hcdf36a7218648e4a471faa36bcb7d8ff690f7b8072efa55158d5414b26704f09;
defparam bigblock17.INIT_2E = 256'h3d3ae9250c1065514d09603137c6174eee29aa5434fff39cc3bf8fe5ec6e3fed;
defparam bigblock17.INIT_2F = 256'h0366ff807274fffb9caf0249deaa8d314cd30e09d7131ace66aa0e97361b715e;
defparam bigblock17.INIT_30 = 256'hb13da69ba52068b18b6de87facf86ae76173900d2162db571e622f98b9e740da;
defparam bigblock17.INIT_31 = 256'ha6a33654055d99215c052b69b3d68914f6ad07ff588084f0a63ad15e4807d7fd;
defparam bigblock17.INIT_32 = 256'he6f3b1eb66429a242ac2b272ccf1b36d4347400244809200036c898a0c32e250;
defparam bigblock17.INIT_33 = 256'h7f7288b3ec4b73c05f2f2431030aeba440b4d008f46b24d6dcc2f68c11a8ffe5;
defparam bigblock17.INIT_34 = 256'hfffb6fd62ff92fff434be8ff5c97fce1e8d4084ed96ec673a4cf01a9c789effe;
defparam bigblock17.INIT_35 = 256'hbfb5da0c544003ecc6a55a8dfff0ffffffffffffffffffffffffffff9fff387c;
defparam bigblock17.INIT_36 = 256'h498d0bb27ad9895d001b01008834413839bff12335f9a681ae04e2468eeba5b8;
defparam bigblock17.INIT_37 = 256'h2d3ea533c7459699666fdbd763e25c532d436ad56ebb0b4c95a2313b83751a8b;
defparam bigblock17.INIT_38 = 256'h4eb891e2ba163833193ccd3e3527e09beb858d8fe8b9759f24a5763a5a2ae1fd;
defparam bigblock17.INIT_39 = 256'h3c60d1eb3259031aff807274fffb3f9c5169b6df4576b73004f406a1f040e2ff;
defparam bigblock17.INIT_3A = 256'h08bc7f9482cc99ec9f141d10d8f3092c2079b4fe6647893b664e2d05bb372042;
defparam bigblock17.INIT_3B = 256'h7b9dd0bda2907b721923739d42eeff100381ca91942e6a1eb71c06015828bb91;
defparam bigblock17.INIT_3C = 256'h0544daa1d4d0e043513d40e518d6f29149d9c9f71a9339a999e15bdba0007e0c;
defparam bigblock17.INIT_3D = 256'h91fc2ba1d490727a3bdc8ba56395298926ea46b7ba89c4d496da585865de0d43;
defparam bigblock17.INIT_3E = 256'hfbaf015ba7d5661fe0c9ccf16d6a68217734316f35954313638f61f03f1fb596;
defparam bigblock17.INIT_3F = 256'hffffffffffffffffffffffffffffffffffff2cbfef956fde3383f442d33fa1a3;
defparam bigblock18.INIT_00 = 256'hcbe14c4e38916500d24a62d951789f54c6bb92468d1ca81ce391fc16ffffffff;
defparam bigblock18.INIT_01 = 256'h097116d64d528dcd6cc98810f8099f17b7b8f438c24e52920fd30011c0805484;
defparam bigblock18.INIT_02 = 256'hc310a459c7ae210ffd647ee7834157902bd0b756e2f03010af36c26922c559b6;
defparam bigblock18.INIT_03 = 256'h1988db3320425530b9e940d90354ff807274fffb37ffd3e6047f7fc33ce66d75;
defparam bigblock18.INIT_04 = 256'h371b0041fb05efeb2fffdfffffa0e2fe2921cc640aec2078acfe66c7a921360d;
defparam bigblock18.INIT_05 = 256'h124000400c1536640602e7bdd412d4948ec99902e2210629f8d44f3806a16945;
defparam bigblock18.INIT_06 = 256'hcb10708af5f0f475e7118ed25895b96e06ba9924873afd1eae82c649babcbcc6;
defparam bigblock18.INIT_07 = 256'h44eb3ebd512ff50703ebc6a4052a38128ccbdb2690ca904e1401d53011c54f94;
defparam bigblock18.INIT_08 = 256'h8b7ffe9f340befeafee72dfbfa935d7f1125eaf4e21fd4899cef82d4c0c497f9;
defparam bigblock18.INIT_09 = 256'habb9c1de3fb9b21c0f9eeb815b9a8a68deb422360ddf49eb291bff02ffffffff;
defparam bigblock18.INIT_0A = 256'h42a95791e67c42d1dafc0d42ae5b8e7200558000a5408f8384df3ac27d3ac9a4;
defparam bigblock18.INIT_0B = 256'h442c4c50a8c8269e53ea386cdea9e1099e9cf8b78460044c4a7f620fa3175939;
defparam bigblock18.INIT_0C = 256'ha95f54c05f7f24c8eb30e56f3c9980e799696b406de60114a449b34f63328d17;
defparam bigblock18.INIT_0D = 256'h6667b1771c0a192adb331dc255c889ed4f59040eff807074fffb9b7b44d2f529;
defparam bigblock18.INIT_0E = 256'h93b6c905a2fcb4ff8cf16d4449233d007f5ae9c3ff3d9560dc960b2c4080a855;
defparam bigblock18.INIT_0F = 256'h16f57bad6ca410010a002f0c2c9089db3b19815fa5168736bba3a2e31aabfd3e;
defparam bigblock18.INIT_10 = 256'h4ccb7dd579ab6378d41a25f9e2ac6b59ae79e78adbda8d89d57c7c4839c86161;
defparam bigblock18.INIT_11 = 256'h02423427a8c732ebebb57412a38037eee8e66aace166dc2e6b3cbadff75a0951;
defparam bigblock18.INIT_12 = 256'h62ef90a252f506ad08189944ac43b86ca1a49f7294cd32bd82a6f48a2eb7e81b;
defparam bigblock18.INIT_13 = 256'h7c93b3699d1959be02512b43001383c1fec000ff95b0fbe7bfc757b5c554fa1e;
defparam bigblock18.INIT_14 = 256'h8ad4b70c2403c41d9717382d000208005124402ad50495745e9ab832e7a0a07b;
defparam bigblock18.INIT_15 = 256'haa105222839956eaf1eea951040961db08be8833e15edf97f364b26e538dba22;
defparam bigblock18.INIT_16 = 256'hfffffe5329f5799773fb5c62279a34ca166607c0f22dd0601f19f0342c539369;
defparam bigblock18.INIT_17 = 256'h6c0c928bacc007b125610c45caa0033c42db1026e86d58294849800374fffb72;
defparam bigblock18.INIT_18 = 256'h1fbb3a53319eebb1c0c0f088e5b87c67a6d7838db200f4aeff5b4dfa90eaf4a9;
defparam bigblock18.INIT_19 = 256'he1f76c0cd608d5e4a95a02e821c01f5e8b12f88480d3e64746f4c126d512a246;
defparam bigblock18.INIT_1A = 256'h8d4b2e543ba12945a80efd617c293e03f0f740e56461be35f8e1ddef8fcfc0f0;
defparam bigblock18.INIT_1B = 256'h88556d519bf73116de4443ae496928c1b480ce2b5c7c14ad80acf571f1b205b4;
defparam bigblock18.INIT_1C = 256'h91b416dc1d0400c06a7ff50cb69319be189a57639faaf21337a70256d4e29f37;
defparam bigblock18.INIT_1D = 256'h3200894901429c0a228da62662fabba1799484d685a204218be43ac5460e9108;
defparam bigblock18.INIT_1E = 256'hdead85bbb528ba4b8129484a604423b2011293a56507a901602101d32a810000;
defparam bigblock18.INIT_1F = 256'h7193eba1ba665ab54609331e7b966aab14faaf1b93c967ab68d8f1e04752b814;
defparam bigblock18.INIT_20 = 256'h800374fffb72b6ffafd0ed0fdd2910d0b8142579d7dd01128b8f22241b7dfa6a;
defparam bigblock18.INIT_21 = 256'hdf4f084dc6ae6c9c960b5200263d23650af9e7282619a2dbb823ed2e5941a957;
defparam bigblock18.INIT_22 = 256'hc085246891c9715bc3006b8271999894d72ea3c1eb3c91738a19e34f623fe262;
defparam bigblock18.INIT_23 = 256'h7b04eb8490d2dc37a4914419000001197d950620943dc8f55d61b06248c36afb;
defparam bigblock18.INIT_24 = 256'h6ad3adb33292069510b52ed4b7ab8f79f168a248c56097fb3a85ec4a44f568ce;
defparam bigblock18.INIT_25 = 256'hecd95f945469d61b9c9e7e908dd8802b874253785c38f9af8d37fbb8b311f875;
defparam bigblock18.INIT_26 = 256'ha1c3963fe392584858c0d8fdb10bc2a16ac66919f63a013c1602ffaef54ad4d0;
defparam bigblock18.INIT_27 = 256'hbabcbe3b049f8f658da017c53c936850b91b0371c451ff255fca287cebca075f;
defparam bigblock18.INIT_28 = 256'hdd58419a4bdea736531d76af63331786a8cb407022e307af020000100005174a;
defparam bigblock18.INIT_29 = 256'h799075d4113900916ba55f72110e903a5ec252c8c4156a81973d7b10d7a8080f;
defparam bigblock18.INIT_2A = 256'h8f545b494050800374fffb72dbff1fb733fa59d3546d9df4ffc8d4ac0797a34b;
defparam bigblock18.INIT_2B = 256'hca00efffd494ff7b89cd66182da86306136044bd256d0edd272a6d0d62dba824;
defparam bigblock18.INIT_2C = 256'hef5e3404cc8eda52267b0d5e1674a8d3c85fe3241c460fd7da36723680002804;
defparam bigblock18.INIT_2D = 256'h22a992ef2baf3484eecacd5d29146821939455dbdb4c0002000102032023a5b5;
defparam bigblock18.INIT_2E = 256'h458aaea491f7b3a49da2904734ede5ada8001577d807ebf1fd30a07c1ec42791;
defparam bigblock18.INIT_2F = 256'h7ffef51fd49fada95fef46a60de559a290d062244c9069e5bf9589c75e1fbea4;
defparam bigblock18.INIT_30 = 256'hbe0e746793d6ef083f655e5f694cc8db0001c180ec0fcf76f4bf59e83fd5a77d;
defparam bigblock18.INIT_31 = 256'h85168515f2393656800500000d0088f0ef40405af44c098f8b12a75be979e5a6;
defparam bigblock18.INIT_32 = 256'hd6187765c3cfa70bdfaa304a34839438e9b315de4dce1312bcfe287114754ad5;
defparam bigblock18.INIT_33 = 256'h673ca45743207903a8358f9eb6208aa0fd2760f06a3e7060088a8fe53abedcf7;
defparam bigblock18.INIT_34 = 256'h4a30416b7818ef3cda41d24e800374fcfb709bffb31d9a7335538cdf7a09b13b;
defparam bigblock18.INIT_35 = 256'h86ebbeae22247fcc4bd975f38cbf28f2f4896d34978bed0087a43b694b152360;
defparam bigblock18.INIT_36 = 256'h5b457476c5ff27d5e971f3d75228644e62d111a6779d6db400dc000000c07509;
defparam bigblock18.INIT_37 = 256'h73cb15505e77b06a1ce3a19c946df91b109c200080002150c2b390af10f8de7f;
defparam bigblock18.INIT_38 = 256'h7e092140b258899b4541c599de0b0d4719b81539d6162e04cc7db71487991a33;
defparam bigblock18.INIT_39 = 256'hf388cda1a2fe4b6e6aba2b331f9cacd59be84e0bda9a57c96299773de2513dde;
defparam bigblock18.INIT_3A = 256'hdb4ce695cf5dd7d2a43cb44d9dcd6d91352300007850d951ea3bfc8ff51fbfea;
defparam bigblock18.INIT_3B = 256'hd856e751941c1caaeacb0034000020020e040507376b3d54103d08601d3ef72f;
defparam bigblock18.INIT_3C = 256'h3e2b5dc3966ebfacfa87ff04a7fa0492421af9e9b0a159a4910c729d5049c903;
defparam bigblock18.INIT_3D = 256'hdd7d02ffd3e59a8651113d561fa076451c0658ac5a6fbc7c5848c4d1ebb35cf4;
defparam bigblock18.INIT_3E = 256'h658c913d4a4d3d25bb2a25426bf049eb4ed9033afe807274fffb1dfe7f54f55e;
defparam bigblock18.INIT_3F = 256'h8e6a0f93236d0037480083bcbdf9e8df97ffd7ffbf959561b4f40aec8098314d;
defparam bigblock19.INIT_00 = 256'h14c00a005b80c511064f8aad632b83831d41cf1de1c842b9c7f4768198b98098;
defparam bigblock19.INIT_01 = 256'h54cbf3995460954799e58e974a7e450d823382507f228d47953eb91f504825b8;
defparam bigblock19.INIT_02 = 256'hdb70b2bf82a3f10accfffcc41b557245e88d7ab7e158d9880c40510e8aad3d69;
defparam bigblock19.INIT_03 = 256'hff82f6cd51001be8fa0e1febf303cabfea046fdbe94ecb3ea8510f95980b373a;
defparam bigblock19.INIT_04 = 256'h00a5ea8bb9d5925d9650a81a89dc2350d4da8913c24d1a0c72470000f8004715;
defparam bigblock19.INIT_05 = 256'h35b6fb0524417076f4582a61aa75f94d5150a00000000d61d351f1c7319837cd;
defparam bigblock19.INIT_06 = 256'h1a8f1160bb0bb1565ef19964478a75b64d114ce72dcaa04a4a0de3ca5f4918f1;
defparam bigblock19.INIT_07 = 256'h477fd3f3479bde8c15fe2aa2156da723416190067245bcc744b1c0700dd57d64;
defparam bigblock19.INIT_08 = 256'h8aecc0959c5a65875977580c3d65db2a24426d3061eb47d90315fa007274fffb;
defparam bigblock19.INIT_09 = 256'h7078422a398894ee08d88a5d8ad98a878db6005bbd41c7e789b02ceeac39a8f4;
defparam bigblock19.INIT_0A = 256'h7d352dc92922477c13370731004011d3588232db586312cf403213332d533398;
defparam bigblock19.INIT_0B = 256'hb6e7bf5f75ebb9484c8ddebfe378af8c313da0dacf75d9eb415238b9e59c8653;
defparam bigblock19.INIT_0C = 256'h8c13db40d39eca9450efb9204425c8973e6bd40da1011fe6f376a9f58783b82a;
defparam bigblock19.INIT_0D = 256'h0009004006fea22af5b3e82b22fa7a9cb6bb083461c1ca379d473f10b7a039ab;
defparam bigblock19.INIT_0E = 256'h2c89d819a8aff7f6767915c25dce3ba179b760aeb7babe8ebab43d9b4f9ac6e3;
defparam bigblock19.INIT_0F = 256'h34d053859add6588b3a01ea216d70f6ca88e1838664ca26996246866452a2025;
defparam bigblock19.INIT_10 = 256'h528c3332b655e4179c0dc1fad34c9a1f186380e275ac164a518b51a182897658;
defparam bigblock19.INIT_11 = 256'hfd807274fffbf51c3bd73d2efb20aabb3624bc4eadfd0a1347c5cb4fbe240540;
defparam bigblock19.INIT_12 = 256'h171ab4204cf40b6c8096c1526327e5051e0b3d2ddb1a26e215c0b30b4858033c;
defparam bigblock19.INIT_13 = 256'hf8947ad454d3b02d48f224a524be03eb248d04a99902f28225bfffa32a67bfaf;
defparam bigblock19.INIT_14 = 256'h68dd5a58dbd72544ada611da995a0521010120c000102631dff4e5376fef6802;
defparam bigblock19.INIT_15 = 256'hc7e1de5fde37aafbec290821da11e66d6ac2f8b70b397015eeb96a23e9064bd1;
defparam bigblock19.INIT_16 = 256'hcea7d6e66abfeb346fff9945d6da27a9db2365f028323e7316a4ac9e5bbf6e8f;
defparam bigblock19.INIT_17 = 256'hb8a1b6604aba3525e2b40549e4894136ff00ffff7fff37f47674fa676dfaffce;
defparam bigblock19.INIT_18 = 256'ha15661d8fad374a6304700a1a560f0197da0956d86ae0da20e9eb9e469262a37;
defparam bigblock19.INIT_19 = 256'hd2b34ae75cf798bbfaaa1248dd49ad6f44b186a2606946f574a5a8c99e36df2d;
defparam bigblock19.INIT_1A = 256'h7e8e9d310d169a3c122616c45ebf301d0809d4a5cfddd6276f5fba443e84e7b5;
defparam bigblock19.INIT_1B = 256'h29eb48d9034fff007074fffb3185b7e6731f3a15fa1a1ea9c24aff9a11673a07;
defparam bigblock19.INIT_1C = 256'hf0d74d2f3476ff33ac109cb10b6ca87cb4f364a40975820d31a8db2a22e23f18;
defparam bigblock19.INIT_1D = 256'he31a6a82b5c5c620bb82b42ff85a35184acb90261b8f8b9d050d49a682dc66a5;
defparam bigblock19.INIT_1E = 256'h4015b3d2671266b6465696f611c31067562b197e6b2b2347300000004075c2c1;
defparam bigblock19.INIT_1F = 256'hbd8c112e0860120b972ae2de10d3f413a8b04a97208bb76f81b280b83440be0e;
defparam bigblock19.INIT_20 = 256'h7fcf8d9eee4073b1c7f37a87fec0fb9f97a8cd2107ee70a79d4ca802e506a36b;
defparam bigblock19.INIT_21 = 256'hd2ca78c42c68349003515f4ed673655d83e8efbf5ff5ed74afffb5dd93f3eadc;
defparam bigblock19.INIT_22 = 256'he490012200000900f248175ffc6a835c540094de5cca2370af26a12e98e5c875;
defparam bigblock19.INIT_23 = 256'h552b0e4c33cc3096fb552752d1a1648cbf2701342537a95ea344fb98ff9bb492;
defparam bigblock19.INIT_24 = 256'hc1ea1e086d93b1958ae2bd5d10e2117eef0f39d2f56e06376a0fe2dcec6c1bd3;
defparam bigblock19.INIT_25 = 256'h172502db40248f6cd8d1284f800374fffb72b2ff210b1bb017cfbc49ca7442c7;
defparam bigblock19.INIT_26 = 256'h69a72fb669101240217a7f9fed104076b7966c4c878bf360263c3f620d65ac4c;
defparam bigblock19.INIT_27 = 256'h55424315b1de3f578f13b243fbff2ffa0a3653c6db9c463e8342356275dcfb50;
defparam bigblock19.INIT_28 = 256'hfffbe9ffffffbff7ffbeebffe99db4599b66ffd5dbffffacf9ffcebfad965994;
defparam bigblock19.INIT_29 = 256'h6b11511433156c5275d92e4f9ae0652842f4226effff3fffa060c0aaebac6fff;
defparam bigblock19.INIT_2A = 256'h5106f3d5fcd44ad41bad7054556ce39a9f79a48899d34b0d89b40e523a5d624d;
defparam bigblock19.INIT_2B = 256'h8ad5403de4fc8fe397bc903942086067e595133197a300006a00109132753db7;
defparam bigblock19.INIT_2C = 256'hd4f17311695dd5558e813284464b324c753856462445c974f05ca07cacc89559;
defparam bigblock19.INIT_2D = 256'h8b0a4a08132464c34b55c759a46430279290bc9cb09717669470a3541a6c4531;
defparam bigblock19.INIT_2E = 256'ha06ba71f939f06bd4429d8495229fcbc2d7bf979bc37fe64eeffc52809e85c55;
defparam bigblock19.INIT_2F = 256'h855e154d2c00f3a642ca08233d6057c58f50800374fffb72d4ffffff0fffe8fc;
defparam bigblock19.INIT_30 = 256'hdd4c4a051aade3fd113143d4f8f79afefbf514bc00c61ef02bcbfe0f80005997;
defparam bigblock19.INIT_31 = 256'h6a6e6ce63c5b4f47000b83004ac9ab73c6240dbec6234b45b73459ace74ec601;
defparam bigblock19.INIT_32 = 256'h7dde82c804c4165a0710863a238dc58966b59f238a3adba0fd9de4dc6152ff6b;
defparam bigblock19.INIT_33 = 256'hab4a2f38c6eca50af0b4815b9323889279d56d194c0e72eaded18deece6268fa;
defparam bigblock19.INIT_34 = 256'h659b6526994a9dfbdfb643bc719c279fe4c91b71e250e9301ab5acbdf09759ab;
defparam bigblock19.INIT_35 = 256'h516db295d8e0ea4dd85d397aff04800fb658abe29298c69075825969ce280277;
defparam bigblock19.INIT_36 = 256'h225a3872e0057a486b652400ad5bb6ce4f0460e73e34de0ec437cf69e6666a9e;
defparam bigblock19.INIT_37 = 256'ha997d43e682ed114a101154fd623403867be53bf5bbab4bd8c4384018234faa1;
defparam bigblock19.INIT_38 = 256'hfa01755f516654784f8338266263503b7e6875f40b7f8b98876000d9465a283a;
defparam bigblock19.INIT_39 = 256'h920c0020dd8611644f8d240022c663ab002e6520d916d640000374cbfb726dff;
defparam bigblock19.INIT_3A = 256'ha9390964fb8eb1223ff06db74b6b5db30059dfaff3fffeb707db012c8c806c8b;
defparam bigblock19.INIT_3B = 256'h026b4f1624df49e8b9019eb23b3aef2047737d16674f6f87bf5dd32f0486e796;
defparam bigblock19.INIT_3C = 256'h182331288279034a2eed58f5632dc1ec1b5c5a1528e7a5923be9b69b3f8e8dea;
defparam bigblock19.INIT_3D = 256'h091e7066cd4afcd45ee8b595d824fd91973320a487325e5db2e69c6ba1fbb412;
defparam bigblock19.INIT_3E = 256'h4013445f0dc2b7d8236db5e7c665ab062c3b7f1b528bb4d961650fb1b9e9e48a;
defparam bigblock19.INIT_3F = 256'h43363cbfd1257668b6ecfb0a29fe48d634eb8f558bb469b5f2e41db1d26f08cc;
defparam bigblock1A.INIT_00 = 256'h6ca41546271475bbe545097406c86f424d0ef1bdff91d6c3a140c1f9d9a448dc;
defparam bigblock1A.INIT_01 = 256'h97222359d88bfe17ca42023d0dc14d09b33e991511fafbac73c87d5cb6f9ac53;
defparam bigblock1A.INIT_02 = 256'h74b1fb70dbff91b659645c52f5001f81850bd1a7d01defa32aa6f373334c7e7f;
defparam bigblock1A.INIT_03 = 256'h293e2199efb490086be0a618fd7d4becc390ed0ca2fb5a23281bdf69a81e0002;
defparam bigblock1A.INIT_04 = 256'hde9b5b8dee11e7987fd438d688c3f298097724abcfd0611b1a58f7020506e181;
defparam bigblock1A.INIT_05 = 256'h630e9471315cd1abe7dcf1d234c0046ad9e42ab302f4a759a3101eb89d146c00;
defparam bigblock1A.INIT_06 = 256'hb83c4ac4e45de0a53181d2ebe363cc756d42b8e0956623af532edc95d5eba118;
defparam bigblock1A.INIT_07 = 256'h101a760e6c9cc6dbfc8d9022d6444a17e8e097dac5d4286b14624a1b190becfc;
defparam bigblock1A.INIT_08 = 256'h902935b822930c26745b88eefeeaa6558a826d995333144b70e398e0ba26bb41;
defparam bigblock1A.INIT_09 = 256'h59271205d4424e6a7a3ac10d8b0bdb65ad56412f8ad94d90a679506702cece71;
defparam bigblock1A.INIT_0A = 256'h02263a2802a874b186acc1f533a401493983a139c788b47045878bad7188b532;
defparam bigblock1A.INIT_0B = 256'h7ac1d593c1e39f4db6d39c29003681091409628c4cb9a62624bd5c4f96a1f52a;
defparam bigblock1A.INIT_0C = 256'he923535f02f1bd807274fffb4a83d615d5f2a458a07071c0b189de222285cbe6;
defparam bigblock1A.INIT_0D = 256'h052904da952904c49518f42090ef6098047e7fa4f8ff244a04430bfd24031658;
defparam bigblock1A.INIT_0E = 256'h64a0f0c20fc3503ebd5a185cb4ee198aa73edf8e09a9a496408bfd60f6aaa16d;
defparam bigblock1A.INIT_0F = 256'hff19912c8e64655ddf20b6a4ffae9c589bfa8306081abe3bb782ccf82e95c5f1;
defparam bigblock1A.INIT_10 = 256'h1fc63c266cf9a6db5d70c3da7fe3df9ded19fdad08bb4fef6fc0f8cfbbd528b3;
defparam bigblock1A.INIT_11 = 256'hd0007126caea8ea53d84d1b7feeb723b2958f8cc489e0c851822c7eac373603d;
defparam bigblock1A.INIT_12 = 256'h2ae303b1986159b1748816f6e3f292f54dfc8e0dac1d8bc2ace2d86cc57b2a72;
defparam bigblock1A.INIT_13 = 256'h502918b34eb13050bba899f94679e5960bf80d6661c432e9eb5288ad314c2748;
defparam bigblock1A.INIT_14 = 256'h87efb0a9ff85d4ff4c78a47f908628e1a28c3358ab859ae8ae43f5c4a5e50d30;
defparam bigblock1A.INIT_15 = 256'hf28d810440e3942909a7ad8a3f461b7615d9b4ad3dfd24c7c806ea6e42733d9c;
defparam bigblock1A.INIT_16 = 256'hdbdd244231e0e8c9185e02b9c8807274fffb560695cbb052cb6a804ec45cabcf;
defparam bigblock1A.INIT_17 = 256'hd383d18168a348297fcf75ae64c30c9968130aef0893206f7ba67c87440b0c28;
defparam bigblock1A.INIT_18 = 256'hb340d3cc9628110e6c7769dac8852f783eeb60fbe5cca634c36da9e4b3cf94c9;
defparam bigblock1A.INIT_19 = 256'h11a3a860b8ed1b6d0e4748d2cb72685caf14fcb05b590513334ab825b40a9d42;
defparam bigblock1A.INIT_1A = 256'h2926428a0b25f4124b8de47b28ab3a392604095c5332af71d058e92f674526f5;
defparam bigblock1A.INIT_1B = 256'h5058acebe359eda99f5bb0c6ad944d442212e1b978b1a43fd9f51760a9485004;
defparam bigblock1A.INIT_1C = 256'hb9684866f0e5fa44397beecd68cd43e92d620e21eec8648711035feb1902f505;
defparam bigblock1A.INIT_1D = 256'hb8dbca723122c7d0cb9a85c8bb3b9ed831c4de9189c511650c72c8de291877cf;
defparam bigblock1A.INIT_1E = 256'hdcd2770a7ea5d273a81b6cf61629be771e7c489b5fd960ab2b83466269c06da7;
defparam bigblock1A.INIT_1F = 256'hacdf7d53c0ac726eff5e57e0d411cbe843c5c5554864fb3457ef939eb64046f5;
defparam bigblock1A.INIT_20 = 256'hfcbd260a04c22be920e41b286989346002e7d5807274fffbe5ffb07533dcd6bf;
defparam bigblock1A.INIT_21 = 256'h3a3468af1ded5ab906cbcb55210c0057d55292398db2b46290f1c0a1a0747da4;
defparam bigblock1A.INIT_22 = 256'ha450fbbd7effff4b950821dd9dcb474333a752c73ab4fa7a8590936cdcb2cad4;
defparam bigblock1A.INIT_23 = 256'hd0003fd542774987d6ac38370751288004c6b419b6d75c6d52c7189c2b447790;
defparam bigblock1A.INIT_24 = 256'h636980c35537976eca9b19710017651c444566838743a0731d5b0125cb4d1a5f;
defparam bigblock1A.INIT_25 = 256'h95443f4cc16f0907d6dc57613d5f45015af11c2aab790ad52ce61829b8aec3a5;
defparam bigblock1A.INIT_26 = 256'he26b8f48fcf0c5b450df6de1ffdae1be1574faa178e785a29c7a3eaaa53f7b18;
defparam bigblock1A.INIT_27 = 256'hdaab7b26a45a9d0053f56db4c9db43756b442b4e16eca5b62687a5a49c401678;
defparam bigblock1A.INIT_28 = 256'h59a6282080a545248b411e1602044d8757633cbcb74fbba53b505ec570cbd1e2;
defparam bigblock1A.INIT_29 = 256'hce701bad4f8c6255d40efa6e01d40fd209215a05a12e6b5beded01c445aaa44a;
defparam bigblock1A.INIT_2A = 256'hc89eb0497fa7316da20c08c23bfd24a41d10e928415d02f2e1807074fffb7a11;
defparam bigblock1A.INIT_2B = 256'haa48fbf274672acc7d9dad179cc610f99a31b6bf8e7c528e954d0a18f42490ef;
defparam bigblock1A.INIT_2C = 256'hc2724ca846a26da636dab56f40ade41159e3469cc76c21a95a52c41698693197;
defparam bigblock1A.INIT_2D = 256'h481e0017889808250060e8db2a7ec2ba98b5a6ef4827af7eaed4744cea16352d;
defparam bigblock1A.INIT_2E = 256'h3c85e657f25ffe06ccb4a5e5baae48d96cf493b7355a634f7cbe16802c2b9b6e;
defparam bigblock1A.INIT_2F = 256'hdeb65bb1395ececedbd4c9f272f9d16f916226779b43306f20ed100d6cf6ad65;
defparam bigblock1A.INIT_30 = 256'h6fff19915e0466926b3447faeb3ba9e2ba0944b85094300530d8db9f1996e71e;
defparam bigblock1A.INIT_31 = 256'h590f36a21763a1b1175157b11aebbcd55acc943872a6b664398b9a460b64792c;
defparam bigblock1A.INIT_32 = 256'h0d1aee91e8f44668dd2f345831edcb62123308f1e025c90a6bcd00da09408951;
defparam bigblock1A.INIT_33 = 256'h74e6fb72c1ffcd428bd5de8ae617cf0adaf15bd565f29e9998b68399af44c58d;
defparam bigblock1A.INIT_34 = 256'hc187578aefa88d8d5640a324ff7d0b3ce35e0d18243c2827881de07915430003;
defparam bigblock1A.INIT_35 = 256'h5818b3c55890ce5815bd8e38397388732648ef1a59519160ccdc7442e8fff228;
defparam bigblock1A.INIT_36 = 256'h70e1a38ff91a266a6aa0de3a4d8aa0e087a24a1c7308bfff822a48c81d99b5aa;
defparam bigblock1A.INIT_37 = 256'hefd6ab8d8cb11c9d514a6d53c701a9d52239c5aa800595c89e83221b2d6cf592;
defparam bigblock1A.INIT_38 = 256'ha7159041572ac7dbd982ea555a9b5cdfc2be779df925f3d1e769c26a189999e7;
defparam bigblock1A.INIT_39 = 256'hdf68c4fd3d62e7449deebab165f5acc8559e9321115ac3f2df4102bbcc8d3112;
defparam bigblock1A.INIT_3A = 256'he93e8171383a8eaa50e25daeb620d36d4a98fad4bb2128c66f41c5bf7d01f636;
defparam bigblock1A.INIT_3B = 256'h9833faaa2ac094005729b243ec48728602b8597ba324073fe445f83adf0f48f3;
defparam bigblock1A.INIT_3C = 256'h53d41458329106aa4df9563589364799db9f67a5a0e94d4426360e01da346590;
defparam bigblock1A.INIT_3D = 256'h5ce9263b800374edfb7219ff9de3bf2ca943b83ebeb258d3b8e730f7674f1dc0;
defparam bigblock1A.INIT_3E = 256'hc2b649ff2da6001d308aee64858a750044acd7734c30c5389904641ba0242f34;
defparam bigblock1A.INIT_3F = 256'h67206dcfa4db12ea482cb7199c0651587f258bb90dc9136a63495814f799d4b4;
defparam bigblock1B.INIT_00 = 256'h2eac0881e36b371dfe891a2f9ea9940dd2b6453fb6559434de621280ad3b40e3;
defparam bigblock1B.INIT_01 = 256'h3f238fa0229e6d3102486d0e7c246a07e691df94e6de4f8ca09cae2ff23502e4;
defparam bigblock1B.INIT_02 = 256'h867c836c9b53caa5a24cd32854cddd900874da3db3be1a500ea4dc40e15f3be4;
defparam bigblock1B.INIT_03 = 256'h7d07fff7382ab7afdeb3739cc8351154e868aaf2a7302d67e15d7f437a1ae556;
defparam bigblock1B.INIT_04 = 256'h75d23702238abcf01e72616acede8c89930002ccaad37854275b48218611d818;
defparam bigblock1B.INIT_05 = 256'he3363d4b7ecf167a1621e29b83d91ad194a3c8e0ec920b116c74d38add5ec001;
defparam bigblock1B.INIT_06 = 256'h85e780651a040d544f7596a8b2477d92acaf940fc608f3ffc748f55306b26a1c;
defparam bigblock1B.INIT_07 = 256'h443b90288f2ddd51334b800374f2fb7295ff071f434fa8e9aa9c28f042044b38;
defparam bigblock1B.INIT_08 = 256'hc9a1b481cb94de764105169b91d730a5eea8958a78c0449411750bc16594aa09;
defparam bigblock1B.INIT_09 = 256'h2f9816b51e7a87f047f6fbd9c0938cfbdcf68c098846b8322ee37fff90db0ac9;
defparam bigblock1B.INIT_0A = 256'h16f56b79fe96cae5d6d39042455362385919005d001940012600b28a31c95a05;
defparam bigblock1B.INIT_0B = 256'he6ad81849776a54688f67133a1ff40de17561f4cfab4735ef8908c5f75e58ab4;
defparam bigblock1B.INIT_0C = 256'hd239d2792fcb0f2450b99e46547295b418a11b7b77d6a20dca6596703a07f998;
defparam bigblock1B.INIT_0D = 256'h5dca11ca46992309b4aae08d05f700007f81b9bda8b1490aac2420b51f1f65f6;
defparam bigblock1B.INIT_0E = 256'h2c2511c1a64f66d3029800ac03008d0e21f98c2dfec3d735f509d1cb18c68aa9;
defparam bigblock1B.INIT_0F = 256'hb41a2506d7bee4c097d9217175c98fa8a89246b8d6245ec231fa53bd07a8eac1;
defparam bigblock1B.INIT_10 = 256'hf6bbd25f8f415ea722138b5b61676b8f8167d47935e166add11d435857851628;
defparam bigblock1B.INIT_11 = 256'h0c44a266960c043b402288155cc9f044800274f4fb7010ffc103a7560a253745;
defparam bigblock1B.INIT_12 = 256'h988affed026bb2b4736ea98ff28e7038142c51a723166e5893901600463da573;
defparam bigblock1B.INIT_13 = 256'hae0e477bce597f3b16fdbca5c0605a37f4400212b8d44616620ddac30684f986;
defparam bigblock1B.INIT_14 = 256'hb3ab97c19373032890d3e549a8769596598d142bea6a8ee83d113d80502d61c0;
defparam bigblock1B.INIT_15 = 256'h24a202a9d2e2aed86c99133ff79a6fd73d6290ecd621389f51ccc318c1d1a63e;
defparam bigblock1B.INIT_16 = 256'h4807cddc8c568755bfddcff2877b6dad668fbeb65f7c2ec932925ec6b516f23e;
defparam bigblock1B.INIT_17 = 256'h185e2ce72c9ba842f6b36dbf18db4229891267c05ffcefbbfd6c93df2ca6e85d;
defparam bigblock1B.INIT_18 = 256'h0eae8f1094e2dc0005b642810d24663d4181c18cf7afa14a64a03abbd431e942;
defparam bigblock1B.INIT_19 = 256'h12e98e336352ae4317d2bed6337db7a8904e46be7f1aa4873f97f6067959908c;
defparam bigblock1B.INIT_1A = 256'h4cc26d5d39329b5b53212e487fcda7bfa4e0e797cb1657374309d6cc6f16272a;
defparam bigblock1B.INIT_1B = 256'h009abd166f2570f5264c05259b7922e31e30e1e84bdb0341fb807274fffb9e5b;
defparam bigblock1B.INIT_1C = 256'h659e36db1a67a0227009aefa96a1735bdb4cb8263557ba0ed3d02da1d8610e6d;
defparam bigblock1B.INIT_1D = 256'h0e45258fd13f0fa9ea58ad5b042bab41b8dc1af6be13fbd43c20154710b76a0c;
defparam bigblock1B.INIT_1E = 256'h98feabe759df7f9f5c82a238ff5c8475567b0ca81cf9e38806a8a00069281a00;
defparam bigblock1B.INIT_1F = 256'h9cf9aa9da185b8aece2714009e33edbd168167d57f839f8e54d8b8eb65636a9f;
defparam bigblock1B.INIT_20 = 256'h35b91841ceb7b3668bceba765cd14b5eae7b98a35cdf64bd8fc92cdaf5945fb5;
defparam bigblock1B.INIT_21 = 256'h48b4a4cb2de048a856db506dc297f86bd7a90ad4fd905efbafdd79e76f6b089c;
defparam bigblock1B.INIT_22 = 256'h089734939024e818ef8cd2f6a961d5bc8c76b099aae2348346cc14df0fdfa506;
defparam bigblock1B.INIT_23 = 256'hf9f838ef7ead2a77e604ad53308ecd4708f72737ce3b9c5b5a8aec23ad2a1c37;
defparam bigblock1B.INIT_24 = 256'h7274fffbf33f5c8854363907aa24e83a356bd58a9c1dfa155cec3481664873b7;
defparam bigblock1B.INIT_25 = 256'ha621b432106ec0a2ac7675a4e511664b18a29bad262332fa61eb445d036afc00;
defparam bigblock1B.INIT_26 = 256'hffe68bbfa3b8a7af98e486852ce9c677c3a8f2e250811f17a377fb0b72cbe062;
defparam bigblock1B.INIT_27 = 256'h0195f88f85494c42f518d05a35d557e3d4c5a8cfa5a9e0f7271ff356147008d9;
defparam bigblock1B.INIT_28 = 256'hc5674e590b21c98a87c426962c23f92f2f0b60d3b54f89234c3d001998a01292;
defparam bigblock1B.INIT_29 = 256'h53d191dc4546f92b74f25a8fa953f356913996b9ca177f442726cffa0039dd6c;
defparam bigblock1B.INIT_2A = 256'h4117adb3657ddbc8895a48a8e673eea4302b673b49b795a365184ec8cec886a4;
defparam bigblock1B.INIT_2B = 256'h809c0c0c67c926b776e56baf1d460794309c3bf36db78a63ca0c2162e5fba851;
defparam bigblock1B.INIT_2C = 256'h95d4f2a67fffe0106aceb58758fd26742029c8e0194e65243c5fccc9a935ffe0;
defparam bigblock1B.INIT_2D = 256'hc9a0a38322b684900ab83f14d06e7acaa3d24130f16b663eb11513f92a10a794;
defparam bigblock1B.INIT_2E = 256'h43dd039af9807274fffbd6962a24d6aa62ed4315a82dd35e84db4b437b7fadbf;
defparam bigblock1B.INIT_2F = 256'h5303231bb58e08a1a4138eee408f147a75a6b8f72a4b04c7abaa26234caa692f;
defparam bigblock1B.INIT_30 = 256'h71fbb6da238a451494093246e48def4d22721d4520d784eb6aca8ac98a98abf8;
defparam bigblock1B.INIT_31 = 256'had631364a489561af074f0a171bf2048a47fe39cf5027a3674af065161e5e6b9;
defparam bigblock1B.INIT_32 = 256'h1f4d163dade7d2711d8807d67f9775efe0573579a8a9eee48a3128cae8008d3c;
defparam bigblock1B.INIT_33 = 256'ha33ab68d0ef2fbe39739f81d1a929ae93c6e58f16635136ce84de456d2f18d80;
defparam bigblock1B.INIT_34 = 256'h089ca278508a458b8c7fc7393ba8f9dfea43d9ecf5aba7411def54b2e8c56cc8;
defparam bigblock1B.INIT_35 = 256'he1218745723e70141b169be2b22a9ece82f6a6d8ac004401b7de336da0bb1198;
defparam bigblock1B.INIT_36 = 256'hcf5b9699a8b91b3b233df1f77b48c4f64151755026a40a76112d718454467295;
defparam bigblock1B.INIT_37 = 256'h7f915280eadaf26e4b83fe12304cd6bf41e4eda3fdd6342cdfeecab84ad6ce64;
defparam bigblock1B.INIT_38 = 256'h2404154a692b585e0330f7007074fffb13f0f429cea1a5bcfc5ec23b820565de;
defparam bigblock1B.INIT_39 = 256'hcda622411d8f868dff65c8fc95993463106fa09a3d1279a6510f760d18223bcd;
defparam bigblock1B.INIT_3A = 256'hcd382b46840bab0d68f456dbd3d596c4d60080a853c78c7f58f548a21a230048;
defparam bigblock1B.INIT_3B = 256'h17abb5e300006945014af24a51a8e7d613db0f953beac90c7d24a84e3db67e94;
defparam bigblock1B.INIT_3C = 256'hcc0b966d71bb5167f6c496b8f9641edd2d98d6e435d5ba790710ba8868e81cec;
defparam bigblock1B.INIT_3D = 256'hecce2ff4ad70f5b86956a029ae92106ddb173b9c24ec87798f382e553c2845f8;
defparam bigblock1B.INIT_3E = 256'h2f4ff62e6210348ce817b4f316485de9c01020a36306509530dc32ab346be9e6;
defparam bigblock1B.INIT_3F = 256'hc7ff012cdbd8cf2a81a6fd82a8cb5ebbd9f616a9362196d16db425424240e008;
defparam bigblock1C.INIT_00 = 256'h2c6f8e5db656ad00190543657094f151c18302ab012f8e981f52c8589a39d5dc;
defparam bigblock1C.INIT_01 = 256'hf12b089e53f11e98fc4d354e2624fa1885684dc70145580ce23c10bfff8ed20c;
defparam bigblock1C.INIT_02 = 256'h4c61c51adf04441b582a8d2c5ee9054a000374f4fb720bffc322f2546b2bb2d7;
defparam bigblock1C.INIT_03 = 256'he232ddfa8161562ad5b756e097d78dab49de9895149c6f749c907860a7a0137b;
defparam bigblock1C.INIT_04 = 256'h809fd7f8cd5c411c9adfab577a060dd248f768b2c6da024880c145434c048248;
defparam bigblock1C.INIT_05 = 256'h57576a8bc28ced115a6caf4e6c42e2a561410ec102c00e121dc093cf6183dabe;
defparam bigblock1C.INIT_06 = 256'h672e446839ae754e151d817be2c9cd9a3deea77e9843fd354471a6b0a5384a33;
defparam bigblock1C.INIT_07 = 256'h2d22b7123df236c2eda20ccc80218c5271b2d52f3561b1121c6607885e896a95;
defparam bigblock1C.INIT_08 = 256'h764813d227022d6d1eac78a33fff00221400ccc03b0a5aa13f532f7b4047ef17;
defparam bigblock1C.INIT_09 = 256'h9517eaba71d27aab926f402c2281ce57b853ff14f455b14f44609c67141c5ef8;
defparam bigblock1C.INIT_0A = 256'hdf3b1267f6a102e77ef450097a50a177a71511ff5db6cf27808ebd8ef8b82b0b;
defparam bigblock1C.INIT_0B = 256'h1e38a45ca6d2bd0bdf9ad71b793bd0cfdf523cfee6637f04f7bfd6433165f367;
defparam bigblock1C.INIT_0C = 256'h584044a013750b952a28ad05439b18258f455d51533d800374f4fb7250ff1e51;
defparam bigblock1C.INIT_0D = 256'h8308a9d46d13811b0021178cd6ca2976d777009ce347d235a113131caea88b0f;
defparam bigblock1C.INIT_0E = 256'h0000993305d45569844bb1fae9c540201972f7d51682fbb7e6ad93274a8e0d2e;
defparam bigblock1C.INIT_0F = 256'h78aba1fed6e94cf6ee8c0a7ddc604ab3ee5949f6a209548142f5d2f11a42a386;
defparam bigblock1C.INIT_10 = 256'heed0247155a7522b53b38d022a9be043d86a47281ca35477528c7104bbff6d7d;
defparam bigblock1C.INIT_11 = 256'h651a72e6750857f596b6408ad1bdb58152d6a81048eb0b3c8d357bd02a2bbb10;
defparam bigblock1C.INIT_12 = 256'h56cd3277daa19c9aeff891bae3b94a0ec32e6a1fc6db2008c062a31f6592c5a5;
defparam bigblock1C.INIT_13 = 256'he78d4ce3207efe65d49e84432c993007095831014cba561042afd8cf7ce6a01a;
defparam bigblock1C.INIT_14 = 256'h9e32efb963145a558ecc5e931cd389cfdeeeb48a9ee0548c004803adc40135e7;
defparam bigblock1C.INIT_15 = 256'hfb7219ff51d990f96599b9fcc6ed68f9b9ac4ad37f7ecea7c99e6c96078c3e82;
defparam bigblock1C.INIT_16 = 256'h83156d9c900bd600c614df6c4c0425286c0da2bb302488165b312245000374f8;
defparam bigblock1C.INIT_17 = 256'hd5661190e506db391b4a06591082a54031c62f6a1763ca67e147e74571e22830;
defparam bigblock1C.INIT_18 = 256'h9e3a0092009c4588aea4460e2e99070d7f8c3b8a02bca3fc9647380932de25cb;
defparam bigblock1C.INIT_19 = 256'he7fc74657436725378330c6bcf8c14013bc7f47bd45e0a236da37bc86a95e46a;
defparam bigblock1C.INIT_1A = 256'h1c20ad4a50402c2f2441d27bc5251a04dd778ec6011892b2bb05599101a4583d;
defparam bigblock1C.INIT_1B = 256'haf809e8c3d21e9f53e94fd0c6a5febfcede4163d09557d355a3851edf0b3e894;
defparam bigblock1C.INIT_1C = 256'h0bd0dce3e0edd5fc717934b8b435aea5dc2425389634b49ddbbd463600414c04;
defparam bigblock1C.INIT_1D = 256'hb399edcb323ffa8b9f0f9f72a7882aa8b70ac8c8a92484a624019122c4904856;
defparam bigblock1C.INIT_1E = 256'hef9b6f2cb7da90cae0c8d8a6c138ccfca369d1a7e305a997ab4d477961cb56ce;
defparam bigblock1C.INIT_1F = 256'h624b800374fcfb70e8fff30e2e704e9cdb72d7583d7557efbddf24ec9b0fa87b;
defparam bigblock1C.INIT_20 = 256'h974d7904897e70a2ee689b0fd120231c09734c11e3889a2483db88262f45dcd1;
defparam bigblock1C.INIT_21 = 256'h9fd7556e2bf6a89f63c836d81b6d2d030bc0f59014ad5a1270f5105e03cbe581;
defparam bigblock1C.INIT_22 = 256'h2195044f002724b8514e0328e7a69d2838e749fc437675948417bf068bd79e1f;
defparam bigblock1C.INIT_23 = 256'h6f460af305a643380fef38c37c3db2d2785a2839796d3f54ae09ae9a154c410a;
defparam bigblock1C.INIT_24 = 256'heb529d0a69effab820907d293173ad15584a7af2868169a91f2d8e196523b7fe;
defparam bigblock1C.INIT_25 = 256'ha36d59b50445ffafd6e504225656c7839d22877ce66dadd5e40e4c9faea3b232;
defparam bigblock1C.INIT_26 = 256'h6e4c2405c4e4fd1c8d1331944f0a015f86d5a85444cba4ebb8d62f57a83cb2c4;
defparam bigblock1C.INIT_27 = 256'h5594a86e07007cf70ae76b6abd0e6dd94d04690fd0211a68c00088511a092882;
defparam bigblock1C.INIT_28 = 256'hcd7c409927a9d7ab2840a8f92c661b91646bc400f8786b7f197bff521b608c32;
defparam bigblock1C.INIT_29 = 256'h25e3437849864b5c0339fa007274fffb4d3a4700b747391341df6377a79af7a6;
defparam bigblock1C.INIT_2A = 256'h276ffa20fedff9fffeed5f0488b928250e2ec098ac7171a7a0f5580c25458b8d;
defparam bigblock1C.INIT_2B = 256'h3daef6e0d62a58a70e80c4a6dd57198434988c1a20d1695ae8db4c296414d203;
defparam bigblock1C.INIT_2C = 256'ha5612a982471eb196591249000b4114090249349ae55a4d6682a8a1d5fffb6a8;
defparam bigblock1C.INIT_2D = 256'he34681e6a471989db0a47ffecfb7e94f99f3bdd7c9bb90f9f463058ac9b2e9ec;
defparam bigblock1C.INIT_2E = 256'hb24a5af0f1649d33ed462103963f674a04cc243f3153c339d7adcba75652d006;
defparam bigblock1C.INIT_2F = 256'h0c24657aa4ad6b6d0308e9b8711f41f46a42e3d9b045f0ca280acf06f7f26c6f;
defparam bigblock1C.INIT_30 = 256'h8091ec1443502ea224ccebe853cc51c4f0a1756c19e9a83057a4a3a6886c9b19;
defparam bigblock1C.INIT_31 = 256'h90243b9a7b1d3df407dd68f51ce99c13c44e699b8c657b2d2d4001f2801d1144;
defparam bigblock1C.INIT_32 = 256'h54727deafbfe496420c832c95f11ed8546a7d4852d6e57d38b3ccff2fcf46286;
defparam bigblock1C.INIT_33 = 256'h2e0b04e33baa26c417186988445d0330f9007274fffb92018b5c57d8e081f2e7;
defparam bigblock1C.INIT_34 = 256'hd77f97fa33ba8715dcb98ef9a625911a4f6b1a18b45490ee60b09c5c75a48561;
defparam bigblock1C.INIT_35 = 256'h3104ff54ad5f36f7ea11b597f916464e58a6fc5a4206c48b1fd68db58263a0e2;
defparam bigblock1C.INIT_36 = 256'h2794ab12777fec5295d1233562cb3b89ede0b1c9e03458015151cc02ff29b58b;
defparam bigblock1C.INIT_37 = 256'hbd553f42b4ac5e04733c0acb2284a3c24beb2aa336dc188ba97aaa3fc4f52666;
defparam bigblock1C.INIT_38 = 256'h96cb3c5de9ba0ca80a31a465e5e331123082255dd9f5286f8fdd20c9da693071;
defparam bigblock1C.INIT_39 = 256'h430d0643ee0e8c81db6b00d60001418088fe4a74f18f4fbdf76e3d975755e8ce;
defparam bigblock1C.INIT_3A = 256'h22a28081d24cc1741733a199f048f0b80f775dd17ec3af35609979deda2bd484;
defparam bigblock1C.INIT_3B = 256'h44ff789fb08d636362f0fd72aa3b876ca946b3419a6a5e6970942979055064e4;
defparam bigblock1C.INIT_3C = 256'he83b259cbf55a1475ade8879aa981d43eabd6d15212f334837b178c8544f09d8;
defparam bigblock1C.INIT_3D = 256'hac777124c929340b0d251b8a2a241f0851284adc033bf9807274fffb0bfdb7ae;
defparam bigblock1C.INIT_3E = 256'hc0103e828fd9c6db024d40200030a3f4ffbbc13afa776cd499e01c6310ee2091;
defparam bigblock1C.INIT_3F = 256'h0b68a821c79d628a1d0c18fe98a7563978c1c4d7017d2af4d85942d6340822b4;
defparam bigblock1D.INIT_00 = 256'hfa42dffbd52c9fce2d63b0c272266cfacd7fab2e57bb60d0231400c2a301a0fc;
defparam bigblock1D.INIT_01 = 256'heff3ad39242681629d7cf0b093c74181cf16116042a8115cd4252c9f58f446ab;
defparam bigblock1D.INIT_02 = 256'h407294dda75b0b1e010aa66ffc8dbabfeed35e5177fb2ed5f62b4dda5c5c3021;
defparam bigblock1D.INIT_03 = 256'h68ba9a90a004022f67fb3fd22f100629419292f499a26db6264d8a246108a306;
defparam bigblock1D.INIT_04 = 256'h2eae8034b691424fa30e20f600148c4c14950f1019707a20a38afc28dab2a712;
defparam bigblock1D.INIT_05 = 256'h86f6b6d79d22fc4054ef39b4b689dc085af1f50d26ae065c00e1fc14db40dd2a;
defparam bigblock1D.INIT_06 = 256'hfffb83f9b3dc57ddfd167b5ed7f38e21af345cd9b9fe9555efe35550129b8bec;
defparam bigblock1D.INIT_07 = 256'hf49390ed00b3a0576ee4752b880a20e63b7d2aa42e48c988595b0357fa807074;
defparam bigblock1D.INIT_08 = 256'h6db4014b9515a6684bcfafbfffba9dafefffdc4b37e1dddc2ffbf117badd1518;
defparam bigblock1D.INIT_09 = 256'h7dd7e94144f1185fc64847097d9476edf8e1141dbddb82ba26fd96332fd8be63;
defparam bigblock1D.INIT_0A = 256'h624c95c76d49c400d5466d1364842ec1af3ab29c9023995bfa000b7315b4917d;
defparam bigblock1D.INIT_0B = 256'hc7ad255ace64d00e35cfb0c3450322e697578633cc7c570c83a9eababe06e9b8;
defparam bigblock1D.INIT_0C = 256'h1ccad128705eb1299d86d3f851295a9938ef430aaa378f5338a38c47c18c88aa;
defparam bigblock1D.INIT_0D = 256'h5ea62e5f1f4feae8f1fc898625762a745b93ed522f04c3723968f3a267aa5555;
defparam bigblock1D.INIT_0E = 256'haac4bdb346f6f58dbd3dfc7958d65b6bd62be3c3b3cf4ccd9b9555f0ec71d74d;
defparam bigblock1D.INIT_0F = 256'hffacffffb81f4cfad6dfbf6e70ddbffff9ddc0cc69adffceff8ffd5bff5f977b;
defparam bigblock1D.INIT_10 = 256'h1b44000374fafb7290ff4f1cff7c99a828d327d424920e531e61ce22b6a8ab9e;
defparam bigblock1D.INIT_11 = 256'hca50615201a492702e6a9d0e8028548563734d09a37a9d2c241bc82bcc435cd0;
defparam bigblock1D.INIT_12 = 256'h7b64d533484ac304072ac485c9545e8dd2d66ad1a00b21aaac2d01380bf22b1b;
defparam bigblock1D.INIT_13 = 256'h38045b4370b0d0dedff16fa76ab8d7598b302260b88843242032b930dc2814f2;
defparam bigblock1D.INIT_14 = 256'h608b20cd663b13289d35683371d83b12504995c040ce958a6720de622892989e;
defparam bigblock1D.INIT_15 = 256'h6b1374a97ca6e29dbd58eb7a99c963fd96f66c531ba6f92df2d1597c3da1d225;
defparam bigblock1D.INIT_16 = 256'hc9a8c1aeab011e3e263fe16672d8c6f025cdc02ed2310552e5d319d3ccdf2210;
defparam bigblock1D.INIT_17 = 256'h5dab9d8563c8691bc2bcbc3a781bf18a301b1eeef17f6df5061abbea1d4eb169;
defparam bigblock1D.INIT_18 = 256'hdd986c5acf03ad1e7fff597bb893e648f2b729ff0bf7d59a4961e59e89605875;
defparam bigblock1D.INIT_19 = 256'h94cc9da42dda51a7d44f613098cc14fae1f77a9002ac50d57c25fd32ffffc0ff;
defparam bigblock1D.INIT_1A = 256'h004661e05806cd64000574f6fb72aaff8db96665c210493452a8a5a96b2a06ab;
defparam bigblock1D.INIT_1B = 256'h572cb13c35c648ad7b6400191ef02c0b030f8001199791601769bc0002c763cb;
defparam bigblock1D.INIT_1C = 256'h46d01110cd6b19b9ddd504dadd826654f2522a7a90c00405796a7a802119299c;
defparam bigblock1D.INIT_1D = 256'hb87d96e86d5223b8d4baa5668963e9ce4cfbd4191f6faddc0baf865c2478d75a;
defparam bigblock1D.INIT_1E = 256'hf53a877ffed797847a84aff87efdd8342a1cffdf534cdd558e50eaab4c9ebf65;
defparam bigblock1D.INIT_1F = 256'hdf0d820ef0f85f6f8e2048c286a9bae7aff40cea29145e00283f7de75bb18416;
defparam bigblock1D.INIT_20 = 256'h55175f194a02b66261898babb62edd80e2d28b9d22229a8f8424f6d240544407;
defparam bigblock1D.INIT_21 = 256'h96ffffcb04cecc8cb07f4c664e8ed2515042cdb76c4c4d5f738e58ca808cc456;
defparam bigblock1D.INIT_22 = 256'hee0e265c25e824b7416b91b13aab6e6777befd4ab3663596b6cba346e2ba1e7a;
defparam bigblock1D.INIT_23 = 256'h12296db2330a4945bac495411e5c84f5894c7b23afa9bffe95a673012c789d6a;
defparam bigblock1D.INIT_24 = 256'ha000ace2422b0a192560dd4f1f3c00037483fb7257ff511119f677a332ebb92e;
defparam bigblock1D.INIT_25 = 256'h5e533975f6f7315d8151a418f44f3497001b009c6ea45007710044ac33754c5d;
defparam bigblock1D.INIT_26 = 256'h556a5e64bd97192e0d3d94cd2ba26a2ab80acb53d0f1f2957898a5327153a7c8;
defparam bigblock1D.INIT_27 = 256'h3f299aed458fbac4d7bb64d8a90e5f6ed8ef9e5c51509021ccca988cef2a9eab;
defparam bigblock1D.INIT_28 = 256'h5c468d37388ac79f05bd42382caa4a92e22e28a69b03f41e9f7fb49bd84d8aeb;
defparam bigblock1D.INIT_29 = 256'h8dffbd2aa917b4413f4c6904415f2dedf7ccd608885a997a23724b6c8ace1049;
defparam bigblock1D.INIT_2A = 256'ha302cc858ede278dc9b240f4ca74fb4f430f96c3243306e6e2c2d943bb9f21e1;
defparam bigblock1D.INIT_2B = 256'hcd472d530194791fa5fbe915ae53fb313cb98e7f4fdc2beb6725b95a894b0ba6;
defparam bigblock1D.INIT_2C = 256'h383a924a952411a3db940f413df7863bd0a959a8340edb4971b89224b069800e;
defparam bigblock1D.INIT_2D = 256'h4dae120bed6b2caab3b540c7983159ddf6dede073e384bafacf65f57b6276dda;
defparam bigblock1D.INIT_2E = 256'ha4a061794ced6724cc04423b4218851e5d692a4d00037494fb7066ffa766f573;
defparam bigblock1D.INIT_2F = 256'h1a918085cf97f99ecfee43df3bc5f865bcbd83cb7db3d060310def3460887a68;
defparam bigblock1D.INIT_30 = 256'hf70d24893e3658cc72541dffec0de9bb2566ef7d68f1c4eee96a548cce0d2993;
defparam bigblock1D.INIT_31 = 256'h34813db82890a28b7f56958d240a4116ea47affe040748a3b5f38a77b8a7592f;
defparam bigblock1D.INIT_32 = 256'hb56b3e4cc17016258f4bfec5b78973bc5f943d654c0890364dcb660d512a73a4;
defparam bigblock1D.INIT_33 = 256'h629ad9362242fd2aaf79838133ab6ea598c6a2b4ff913b1dfa938bbf325f44fc;
defparam bigblock1D.INIT_34 = 256'hd3bac7d4963dcb989018430a9198a9d26592a3b18a3ff4fab4cc9262232d8cbb;
defparam bigblock1D.INIT_35 = 256'h0521aa412aa9c8891a0c545f13bdf6925f04880cb416e36d69a804885f7c460e;
defparam bigblock1D.INIT_36 = 256'h1f71d012b3d0469fe73218cb23d28be64f72cb5457ebd34bdc49919180c21839;
defparam bigblock1D.INIT_37 = 256'hfffbc6835dad88e871c31b2c3deeff2d13b4580e5792758e8d71c610291303c7;
defparam bigblock1D.INIT_38 = 256'hf43106eec060947c77a4552b2c4c0cafdbbc18411792e9834add0351a0007274;
defparam bigblock1D.INIT_39 = 256'h6b50596f356cd91c92e2df74871875752a75fe44b6bb209867392aabf2ce1990;
defparam bigblock1D.INIT_3A = 256'h3a3ac12c34ad45de6ce031cec57ce504eea9411446db136e8414bb4817d82a1c;
defparam bigblock1D.INIT_3B = 256'h8e459fdceb7404c90c45389d9bd1a5016b031736c71806b1099ec03724203a1a;
defparam bigblock1D.INIT_3C = 256'h385cd4ee14eca1d98821afc85bb72cfd70141d7e587a60cae0585e6b620f1743;
defparam bigblock1D.INIT_3D = 256'h924d3ff25bfff9fdce60d1e111f6f2d9f9fea85bfafbbebaad8eb992921252e6;
defparam bigblock1D.INIT_3E = 256'h587a06e22200b845f491c521344a41f64a6b64a43691139212006d0298bf136d;
defparam bigblock1D.INIT_3F = 256'h48b9b2f1903a27b1227bee9e13e4d7ce7addedbdc5ff55aa872ba35a8770dab5;
defparam bigblock1E.INIT_00 = 256'hffe9fc735912a3048e8cb691313a61cc8c518d668d2a8584a9017a3e70b35974;
defparam bigblock1E.INIT_01 = 256'h032cac807274fffb624b66d0e6cb1db2a1c12e90380832e18a674ea569a9342e;
defparam bigblock1E.INIT_02 = 256'h08bfc11309406813846ee84b2d107343bd0d660c18a33b9d1ac21558e1884cdc;
defparam bigblock1E.INIT_03 = 256'h9b67f9b6813c005d18044809908304652fe35682d1efba2f74c653cec4baffa3;
defparam bigblock1E.INIT_04 = 256'h9e695d679bac58671090959f82546cc7c211162e6c976f7f6f1f381f5670b48d;
defparam bigblock1E.INIT_05 = 256'h2fccfa7affb7c2cb65e74338f94e0cc820a7ac8e0bc72451538b754c85d2c763;
defparam bigblock1E.INIT_06 = 256'hd7a072a87d5287d788803744300d9cc11b9f1cfb429250a1ee86fff9b387e660;
defparam bigblock1E.INIT_07 = 256'h540716f58a7727cd2a170c0b29c80000001995a4a20d80deca97daa4cec3fb80;
defparam bigblock1E.INIT_08 = 256'h60d336f8c6104911c039ed00689e02f5874351c328ceb890a14fde25a7280245;
defparam bigblock1E.INIT_09 = 256'hdd3a7a1a67f4d5c77d75b39d59fe26215aa5d766e421459c3bda90431e95a395;
defparam bigblock1E.INIT_0A = 256'h5137bc4e87db79290efa4a53b6d2098d92f04ed4d43e7a2bffb79676a924b1ca;
defparam bigblock1E.INIT_0B = 256'h1e4849854a5c0302bb007274fffb8041009000006b803348d9dd001874892090;
defparam bigblock1E.INIT_0C = 256'h114a9c18bb380e70d202b0782412876ea05a987471a78963260c04c33b8915e2;
defparam bigblock1E.INIT_0D = 256'h6bfb2a9ca4cd23340c1a18ea50b76e9c42de56949ec6d93a9a2b1bb28724c835;
defparam bigblock1E.INIT_0E = 256'h3bfef827653f418a65b48b43fdd52725d4e7aaf5c3b2d9a1729fb15a5382c468;
defparam bigblock1E.INIT_0F = 256'h73a3a00851358b99b741ab98db690046a2c14735b1f4dca84bc379898612c257;
defparam bigblock1E.INIT_10 = 256'hb596d1df6763956a662948da090b7c652140008180a8ea014d8df493ffacb303;
defparam bigblock1E.INIT_11 = 256'h7eaf426424699efa3e0e9196ff01474e36ad552556a9bb503b33eab72d886179;
defparam bigblock1E.INIT_12 = 256'h7a7da2f65aa8fd6ee46f5b74a857a2da67fbee953904b849498f7a499215aeee;
defparam bigblock1E.INIT_13 = 256'h6012f0115cc02a12945f723b01907a1fd23a05c1d34941c60c24d7f81e579bf6;
defparam bigblock1E.INIT_14 = 256'hfced6baf5134531cf1c5a8d5f172f10bc49f555c8ece6e95b925a291000aa800;
defparam bigblock1E.INIT_15 = 256'h24291b471b62151051e659da0312cd807274fffb132cbccabc103190db667265;
defparam bigblock1E.INIT_16 = 256'h26e0a7f7e47233f3792008029d9d845298911c34876dc066a44d69a718f5724c;
defparam bigblock1E.INIT_17 = 256'hdddaf37f1fdf0df1f083fc781433c103167466c912c373c9393d22ff3353ca61;
defparam bigblock1E.INIT_18 = 256'h01803c2a9ee90700b9df6b535b57cd4f8bdc6b38c14cffa605df907c3e00239e;
defparam bigblock1E.INIT_19 = 256'h220e9e45162548c69a2b8d28592f1b5702c982cb3e09b844b100018101c55000;
defparam bigblock1E.INIT_1A = 256'he2f50ef70b3840c2ee386c0f6c47b44a89c271294d4347a94bc9a0b23160821d;
defparam bigblock1E.INIT_1B = 256'h0c71a2c70ddb1e956b0805d91ac2b1255d74c195c975a6905ea228ed69f37dc9;
defparam bigblock1E.INIT_1C = 256'h0400b7547d73498346dc1ce614d9b64104e8404be50daace12ff3f84d22374d2;
defparam bigblock1E.INIT_1D = 256'hec212efb28bfa7ff766eeb5f7246627134d5b895eb84a359a0ef9ba8463d0007;
defparam bigblock1E.INIT_1E = 256'h747e57bba167add861149aecc8539d78910e3738bd487ed8add2287ea52b8d5d;
defparam bigblock1E.INIT_1F = 256'h71a6810b264c04c7cb8a16e11638512858dc02e5dc807074fffbbf9fa576cbd3;
defparam bigblock1E.INIT_20 = 256'h8fef0acefb39a9bd2da721957ed621f59422ff46911a2c99241607eee8662469;
defparam bigblock1E.INIT_21 = 256'h0001801005011ca631bcb7f2e47342ac0333dad5058c98bca8e48fffa8565087;
defparam bigblock1E.INIT_22 = 256'h415b8cd7eb7d2581028beb312a12e8a1720785dec2921ec0b85674fcc269c7d3;
defparam bigblock1E.INIT_23 = 256'hdd1c0c67ac16a8b6dcd6472061ee9b5cb3b085263a50585c52d48c2ff2ab4969;
defparam bigblock1E.INIT_24 = 256'h31c3ae96d59c472a8c36c7af09438a4d20eced08ea762b25c267bc3e810654ec;
defparam bigblock1E.INIT_25 = 256'h32031197141a265131fadb4905460e80fff8ffffffffffffffff7fff20f46c8f;
defparam bigblock1E.INIT_26 = 256'h5552e717b848791692b8117cfc4944a1000170060f2c8b3a170452ab86550954;
defparam bigblock1E.INIT_27 = 256'h508847c3a70b0236d3e995c8834350ca172396addae216626e5cbeca3cbf950e;
defparam bigblock1E.INIT_28 = 256'h2fff4623814652cc7362bb5b95849176fe3ad86655f55e4b22f7bdff6e48ff9b;
defparam bigblock1E.INIT_29 = 256'had885b085ae8c60c776c4c4526806618021bb819232e5b493943800374eefb72;
defparam bigblock1E.INIT_2A = 256'h07b0c5861039ab2e03fbb501f3be35502dafa9b1d228110977338551499f1498;
defparam bigblock1E.INIT_2B = 256'h958a431e3ebca236181b0a1e000901004472b3b9b0b5df5f8166718ad3e8f28c;
defparam bigblock1E.INIT_2C = 256'h591cf6e2fd42a48616b2ae1de36b352c242869b6cb837035c1dba15ac3be50fe;
defparam bigblock1E.INIT_2D = 256'h35a19a8f94ead5ccb28d427da11ced84b0908ef52c48d3f478291040f838cd3a;
defparam bigblock1E.INIT_2E = 256'h004e33c429cf56ca1ca10eabccc6dc396a85d81f2204e43ac67f65512d4b1aa6;
defparam bigblock1E.INIT_2F = 256'h4716576d064e50000600d9cc2c49cf27c7dd95e24c61190f504964cf752848da;
defparam bigblock1E.INIT_30 = 256'h3f71d38c8d919c5ffdb2b6c1c28de2d0ef1969c3d2d7ae0744714b4238c674ac;
defparam bigblock1E.INIT_31 = 256'h9d6248b30219f0b55cc7662de704f485dbd21ee2d382eb5ac74f1c9bb34bfcae;
defparam bigblock1E.INIT_32 = 256'h000374fdfb722eff75cdf26e8e50d15a5a6aa93c855d0b4475688be8ac9197d7;
defparam bigblock1E.INIT_33 = 256'h2bbf317314986d586b8878a0c6180f6a4c95c2465a24e21b281c86165ac9a53d;
defparam bigblock1E.INIT_34 = 256'h9c9e7b4cc6d37c9900f80b52a69c246d001781b0fd020bbdbf8e6501a9a64d98;
defparam bigblock1E.INIT_35 = 256'h9fd1a1bbbf8a1d46b5ede84501de0126e3c40001014240e88743a1468da65f72;
defparam bigblock1E.INIT_36 = 256'h72d97b96e1143d6451bc031e2435489e2b0f40d2b35d531fabeebee31b1f894b;
defparam bigblock1E.INIT_37 = 256'h31ab2c432a1b65a9ed2edd31c4fc3c0fce69a447b5ae185ef88567efc7966f15;
defparam bigblock1E.INIT_38 = 256'hffff3fff967ada96c79589f2ffe99adf0748abd589faf1a6a8ea6c84e583a979;
defparam bigblock1E.INIT_39 = 256'h614913bb46d7d1655cc9b0be866c7ae70821b9076113b682dc918400ffffffff;
defparam bigblock1E.INIT_3A = 256'h63e7d072c9e60d6e19ee5565a4b120239f973a19248e49260dceaaca80084bc2;
defparam bigblock1E.INIT_3B = 256'hfc591034a9e8a91811e4ac41d16322bebce02fc89a52166515a18aebadae20cc;
defparam bigblock1E.INIT_3C = 256'h89455b396a41800374fffb7242ff72a3a14e419996854db7d6548e230047a974;
defparam bigblock1E.INIT_3D = 256'hbe1df6e16f8fff8239e314a06da87688fe20263c2f6d4e552810670c81db1818;
defparam bigblock1E.INIT_3E = 256'h407c7e6155dccbbca33e64df58c1e115088344f968f038db00114080b33af21e;
defparam bigblock1E.INIT_3F = 256'hbd37b4cbe29a92171dcb4207acc5169146fd138d6603e1b10501400031105c13;
defparam bigblock1F.INIT_00 = 256'hf999d4326ef7dd711ef39c05b6f58eedd0ca67718ee644bd9e49ba979a3c8ff2;
defparam bigblock1F.INIT_01 = 256'hb9105b31b4834184e747fd49b31479d4fd80dc8e22caca45cdd301d10d09dd87;
defparam bigblock1F.INIT_02 = 256'hff02ffffffffffffffffffffffffffffffffffff74ff134f35ea1bd6ffc417ff;
defparam bigblock1F.INIT_03 = 256'h005508003e705b282d80308e97303afee412cc243c3bf722e6a16da046e30000;
defparam bigblock1F.INIT_04 = 256'h160c6e19bd248022fdbec615d31c951baac7f0197b92a578e79240b14e9b33f4;
defparam bigblock1F.INIT_05 = 256'hee7c3fda026bee2133e42153e868356d963fc00e3a2fdb6af0b09b800f7521e9;
defparam bigblock1F.INIT_06 = 256'h5708621b881d8b475ac1d14c800374fffb704fff3a99db04906da1236b382d46;
defparam bigblock1F.INIT_07 = 256'hb3527dbb33f97fc6baa3877a58b6296414b06d687b077a80c6201b6a4bd9c912;
defparam bigblock1F.INIT_08 = 256'h00235a0049c7cce905f33fcacafdd9e082a2338a694ab3dc5ad26d20b7244201;
defparam bigblock1F.INIT_09 = 256'he09e71c382542ba340307a14d7450b06091ecb92e4451dd19812060c8a920000;
defparam bigblock1F.INIT_0A = 256'ha079ea1ed5d557d9dbc86637344a7bc19a6c8aef72d298ffedd19a2aab1dcabb;
defparam bigblock1F.INIT_0B = 256'h90b03488d5d8175eb69a67edd5fc70adb3cf5dd70fb53b165fd7c703775eb7c3;
defparam bigblock1F.INIT_0C = 256'h957beac5e9d0b91b6d2a36e3e00cffffffffffff1d7facd5f7764faaa03c6dc8;
defparam bigblock1F.INIT_0D = 256'h6e5121d9e3b4ca8e7b83596ddd0da22d0000a090c64c3acddca26616f98e8584;
defparam bigblock1F.INIT_0E = 256'haa203b504d6388e9fa8b980c02939a56f0f37a0a5bb697ece4772df0c2b44ae6;
defparam bigblock1F.INIT_0F = 256'h62460ffbe56e0e25fb7e85e3af8a9aa3a3669922b31a45ce8d8dbe96bd69eb59;
defparam bigblock1F.INIT_10 = 256'h6cc61d310e4c05252b6a1c822f98318851db03e0ff807274fffbf6f534f45244;
defparam bigblock1F.INIT_11 = 256'h2db99082f6b48d4e493c7750f4158ab792f05baf3db824289c13896d607220b5;
defparam bigblock1F.INIT_12 = 256'h1a424a1249000602c60196010147a8d628276ea313c6794e030caa0b7d471b4d;
defparam bigblock1F.INIT_13 = 256'hdf589430e506d0a12247d094af7d36ac8297269b01b9660e9901517c8d03c1a3;
defparam bigblock1F.INIT_14 = 256'h6a3d4a22d91573f90bb59f9ac9e37d49c20893143d6154307e436ddb0857eff1;
defparam bigblock1F.INIT_15 = 256'h56a02dad34a0f6df36f39c928824fe942dec3fd4bfdeffc2888bd4affd4891d1;
defparam bigblock1F.INIT_16 = 256'ha820c580ff101f5db233de01975843ce15ca449a3342cb0b8997d35bb510f4ef;
defparam bigblock1F.INIT_17 = 256'hba3182ee3ed8299b63da6ef15cc05bc82d2a2123f0e804d1bd851d5e5517241b;
defparam bigblock1F.INIT_18 = 256'h91c4989813bb87c514077469bb6a239e324abbdf5c7ec8220835a42210b20d0b;
defparam bigblock1F.INIT_19 = 256'h59f488d22eba29956e8963ef99bafeb92cbf74a215cd7457e1afcfaffe64df2c;
defparam bigblock1F.INIT_1A = 256'h886d6069a0be6ac7892f064d05262b571a025d28c92f415a03abff807274fffb;
defparam bigblock1F.INIT_1B = 256'heff576d06ef138b2380d3d9c947eb23600d88388f748099996f5e0bf1a015c81;
defparam bigblock1F.INIT_1C = 256'h121c552e43473c15b08cc8c45e07db3e9ff88b7e1c50620ad58e880856079a6d;
defparam bigblock1F.INIT_1D = 256'h676028b362825f2ae27f313470e3505c2f007252bc5149d4ddd925764014d645;
defparam bigblock1F.INIT_1E = 256'hebcf5335e4dec76ed03be9a2b6c30b81ae72e91c49a9108a953ab50ee2ad6884;
defparam bigblock1F.INIT_1F = 256'hdc7fc9ef3cec9a9aa746ade12d555c661a83c69180e123547b0ed3b79a95e31f;
defparam bigblock1F.INIT_20 = 256'hbfdb9fd75b3545fe272a87280b23b4dc5fd850cb9e8c131c6b6ed3cb472df28a;
defparam bigblock1F.INIT_21 = 256'h7b191daf67732de5672adab9b479729bef0d6398625d51b8bb7a30a5d61733b0;
defparam bigblock1F.INIT_22 = 256'h8d7ece6552fd377bfffec6e76afd5ae5fabffa797dffd4cf79cfbfeeae65fd67;
defparam bigblock1F.INIT_23 = 256'hff807274fffb579c189e8bd2944fc0c98d939e3ce212b585b6da1b6d92497e00;
defparam bigblock1F.INIT_24 = 256'h2a068000ea9090ed00b7c5806fb4611d760d25063b772b042d58c9284bdb02d9;
defparam bigblock1F.INIT_25 = 256'hdad9ade5230a1c6d4f58dceec5f23d891504136c9a508799501e1099325d75d3;
defparam bigblock1F.INIT_26 = 256'h906b18ea817b5b42a5c2b6945a145f0d250a84a18a2d4cd5ee22a112393118e2;
defparam bigblock1F.INIT_27 = 256'hd654518f06e55c171d707876618514435c781ec28b90805739466508eab0cace;
defparam bigblock1F.INIT_28 = 256'h2daba05bf132827e88ce9ec2842e72c486ce37980b39a30eab73e1ec9e712cb2;
defparam bigblock1F.INIT_29 = 256'hd7ae87ad798562df36c9097c1cfcaf376cc65f79e2e53e95245c14fb3386bcae;
defparam bigblock1F.INIT_2A = 256'hb8846cde4689a41a571915e35b6a671e6833b9878d2c9cc3bd2fb9fb3da4696b;
defparam bigblock1F.INIT_2B = 256'h1b6d924986008d65e6cb94a5ffe205f7eecbd24925a1fffe20cf2871d614c7bb;
defparam bigblock1F.INIT_2C = 256'h06fe36661de1a83f29744b92702759d81747d230c18aa168d687ad7a01fcb6db;
defparam bigblock1F.INIT_2D = 256'h066364580637fb007074fffbabe4e5788abc46b7692a257595d4dca245914a81;
defparam bigblock1F.INIT_2E = 256'haba6940d584b31baf0000f1e8f2c010c8780601901910016c7bccb0346030000;
defparam bigblock1F.INIT_2F = 256'h49b09e700d49d2a658d96e13abaf8f89dd5a9d71b68b29c604cad4340422d756;
defparam bigblock1F.INIT_30 = 256'haf5afb7316ca51c9cbe58ff45ff2d7fb2ad67971b043a6eb3155acb49fbcba25;
defparam bigblock1F.INIT_31 = 256'h3fdd5357ab4641a314f1dbe97c9fbf43bdeb54e8ff636c276d4ad0e3ff837f3f;
defparam bigblock1F.INIT_32 = 256'h3295548c4e189052250bd5be1b070c257202936626db8f69c0912437f92134bf;
defparam bigblock1F.INIT_33 = 256'h68a652a9d62bd499f3e69c45db5b5cb2b3f6d1f2eb849eacfae4b94e14aa797b;
defparam bigblock1F.INIT_34 = 256'h91cac3476bec22ef094037a657fdae3c4f96402e3b3561976b5ef678b2bba32b;
defparam bigblock1F.INIT_35 = 256'h325acb27b831f9e682f3cb7f45edfdf0482ffaa24d1699c8cc0d7a1111bdaefc;
defparam bigblock1F.INIT_36 = 256'ha93ea22f40a1f46f2de1d12a7a390ee778392120e6f4b696e47148c0029311ec;
defparam bigblock1F.INIT_37 = 256'hbae1e0eb0a1131205def222c80037485fb7220ff3147d1969249353604613413;
defparam bigblock1F.INIT_38 = 256'h41dddbe7e4f6190ebd5351d2db4438ea0194eef4810d5aa8a6201b774d350000;
defparam bigblock1F.INIT_39 = 256'hab0d9a61ceba77102437139440aa74d4e90f44b19d6d3d0784d3cdfd087bfd32;
defparam bigblock1F.INIT_3A = 256'hac29efff9ff13939fe9d3e9cf87e9f08ba6d369495a7d167d8ec3e97d2734cfe;
defparam bigblock1F.INIT_3B = 256'h6083f7fcafa84eb1acd03b29094436066af7391b185238026a1859b8c51bebd9;
defparam bigblock1F.INIT_3C = 256'ha2a06552ab52461092807182dcf410dcea776282d24ead34928822683fa08a75;
defparam bigblock1F.INIT_3D = 256'h5a252b5dfe9854f5705a1f80ee6aa05af2480a4f57b71245d5f354bc850961aa;
defparam bigblock1F.INIT_3E = 256'hee7d233c1e56ea0b2a8fdac46cf5fabb3e16d2b72a0cb2bdd0f7ff1a17dff230;
defparam bigblock1F.INIT_3F = 256'hcb46e8c13ba888d668a06f0835d19b1226b5d4c6b6931b8d1417a127c47590ba;
// synthesis translate_on
*/
endmodule
