// 
//  MAC_MP3: A Low Energy Implementation of an Audio Decoder
//
//  Copyright (C) 2007 McMaster University
// 
//==============================================================================
// 
// This file is part of MAC_MP3
// 
// MAC_MP3 is distributed in the hope that it will be useful for further research,
// but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY
// or FITNESS FOR A PARTICULAR PURPOSE. MAC_MP3 is free; you can redistribute it
// and/or modify it provided that proper reference is provided to the authors. See
// the documents included in the "doc" folder for further details.
//
//==============================================================================



`timescale 1 ns / 100 ps

//`define DATA_WIDTH 16
//`define ADDRESS_WIDTH 10
`include "defines.v"

module requantizer_coefficient (
	clock,
	mem_en,
	address,
	data_out
);

input clock;
input mem_en;
input [`ADDRESS_WIDTH-1:0] address;
output [`DATA_WIDTH-1:0] data_out;

// Instantiate the RAM
RAMB16_S18 requantizer_coefficient_RAM (
	.DO(data_out),
	.DOP(),
	.ADDR(address),
	.CLK(clock),
	.DI(16'h0),
	.DIP(2'b00),
	.EN(mem_en),
	.SSR(1'b0),
	.WE(1'b0)
);

// Requantizer coefficient
// synthesis attribute INIT_00 of requantizer_coefficient_RAM is "256'h24FF21BE3D2336F330EE2B172572200035902B9D223432CC229E285210000000"
// synthesis attribute INIT_01 of requantizer_coefficient_RAM is "256'h30B12E9C2C8D2A8428802684248D229E20B53DA639F0364A32B42F2D2BB72852"
// synthesis attribute INIT_02 of requantizer_coefficient_RAM is "256'h2A682935280426D625AA24802359223421113FE13DA63B70393F371334ED32CC"
// synthesis attribute INIT_03 of requantizer_coefficient_RAM is "256'h3EAC3D593C093ABA396C382136D83590344B330731C630862F492E0D2CD42B9D"
// synthesis attribute INIT_04 of requantizer_coefficient_RAM is "256'h2A6029A928F3283E278A26D62623257224C02410236122B22204215820AC2000"
// synthesis attribute INIT_05 of requantizer_coefficient_RAM is "256'h3630356D34AC33EB332B326B31AC30EE30312F742EB82DFD2D422C882BCF2B17"
// synthesis attribute INIT_06 of requantizer_coefficient_RAM is "256'h215820F1208B20263F803EB63DEC3D233C5B3B933ACC3A063940387B37B636F3"
// synthesis attribute INIT_07 of requantizer_coefficient_RAM is "256'h27E6277B271026A6263C25D2256824FF2496242D23C4235C22F4228D222521BE"
// synthesis attribute INIT_08 of requantizer_coefficient_RAM is "256'h2EBD2E4E2DDF2D702D012C932C252BB72B492ADC2A6F2A022996292928BD2852"
// synthesis attribute INIT_09 of requantizer_coefficient_RAM is "256'h35D7356334F0347D340A3398332632B4324231D0315F30EE307D300D2F9D2F2D"
// synthesis attribute INIT_0A of requantizer_coefficient_RAM is "256'h3D2E3CB73C403BC93B533ADC3A6639F0397B39063890381B37A7373236BE364A"
// synthesis attribute INIT_0B of requantizer_coefficient_RAM is "256'h2260222321E621A8216B212E20F220B52078203C3FFE3F863F0D3E953E1D3DA6"
// synthesis attribute INIT_0C of requantizer_coefficient_RAM is "256'h2645260525C725882549250A24CC248D244F241123D323952357231922DB229E"
// synthesis attribute INIT_0D of requantizer_coefficient_RAM is "256'h2A432A0229C229812941290128C128802841280127C127812742270226C32684"
// synthesis attribute INIT_0E of requantizer_coefficient_RAM is "256'h2E5A2E182DD62D942D522D102CCF2C8D2C4B2C0A2BC92B882B462B052AC42A84"
// synthesis attribute INIT_0F of requantizer_coefficient_RAM is "256'h32893245320231BE317B313830F530B1306F302C2FE92FA62F642F212EDF2E9C"
// synthesis attribute INIT_10 of requantizer_coefficient_RAM is "256'h36CE36893644360035BB3576353234ED34A93464342033DC33983354331032CC"
// synthesis attribute INIT_11 of requantizer_coefficient_RAM is "256'h3B293AE33A9D3A573A1139CB3985393F38F938B3386E382837E3379E37583713"
// synthesis attribute INIT_12 of requantizer_coefficient_RAM is "256'h3F993F523F0A3EC33E7C3E343DED3DA63D5F3D183CD13C8A3C433BFD3BB63B70"
// synthesis attribute INIT_13 of requantizer_coefficient_RAM is "256'h220F21EB21C621A2217E21592135211120ED20C920A52081205D203920153FE1"
// synthesis attribute INIT_14 of requantizer_coefficient_RAM is "256'h245B2436241123EC23C723A2237D23592334230F22EA22C622A1227D22582234"
// synthesis attribute INIT_15 of requantizer_coefficient_RAM is "256'h26B0268B26652640261A25F525CF25AA2584255F253A251524EF24CA24A52480"
// synthesis attribute INIT_16 of requantizer_coefficient_RAM is "256'h290F28E928C2289C28762850282A280427DE27B92793276D2747272126FC26D6"
// synthesis attribute INIT_17 of requantizer_coefficient_RAM is "256'h2B762B4F2B292B022ADB2AB52A8E2A682A412A1B29F529CE29A82981295B2935"
// synthesis attribute INIT_18 of requantizer_coefficient_RAM is "256'h2DE62DBF2D982D702D492D222CFB2CD42CAD2C862C5F2C382C112BEA2BC42B9D"
// synthesis attribute INIT_19 of requantizer_coefficient_RAM is "256'h305E3037300F2FE72FC02F982F702F492F212EFA2ED22EAB2E832E5C2E352E0D"
// synthesis attribute INIT_1A of requantizer_coefficient_RAM is "256'h32DF32B7328F3266323E321631EE31C6319E3176314E312630FE30D630AE3086"
// synthesis attribute INIT_1B of requantizer_coefficient_RAM is "256'h3568353F351634ED34C5349C3473344B342233FA33D133A93380335833303307"
// synthesis attribute INIT_1C of requantizer_coefficient_RAM is "256'h37F837CF37A5377C3753372A370136D836AF3686365D3634360B35E235B93590"
// synthesis attribute INIT_1D of requantizer_coefficient_RAM is "256'h3A903A663A3C3A1339E939C03996396C3943391938F038C7389D3874384A3821"
// synthesis attribute INIT_1E of requantizer_coefficient_RAM is "256'h3D2F3D053CDB3CB13C873C5D3C333C093BDF3BB53B8B3B613B373B0D3AE33ABA"
// synthesis attribute INIT_1F of requantizer_coefficient_RAM is "256'h3FD63FAB3F813F563F2C3F013ED73EAC3E823E573E2D3E033DD83DAE3D843D59"
// synthesis attribute INIT_20 of requantizer_coefficient_RAM is "256'h2142212D2117210120EC20D720C120AC20962081206B20562041202B20162000"
// synthesis attribute INIT_21 of requantizer_coefficient_RAM is "256'h229C22872271225B22462230221A220421EF21D921C421AE21982183216D2158"
// synthesis attribute INIT_22 of requantizer_coefficient_RAM is "256'h23FA23E423CE23B823A2238D23772361234B2335231F230922F422DE22C822B2"
// synthesis attribute INIT_23 of requantizer_coefficient_RAM is "256'h255B2545252F2519250324ED24D724C024AA2494247E24682452243C24262410"
// synthesis attribute INIT_24 of requantizer_coefficient_RAM is "256'h26C026A92693267D26662650263A2623260D25F725E125CA25B4259E25882572"
// synthesis attribute INIT_25 of requantizer_coefficient_RAM is "256'h2827281127FA27E427CD27B727A0278A2773275D274627302719270326ED26D6"
// synthesis attribute INIT_26 of requantizer_coefficient_RAM is "256'h2992297C2965294E29372921290A28F328DC28C628AF28982882286B2855283E"
// synthesis attribute INIT_27 of requantizer_coefficient_RAM is "256'h2B002AE92AD22ABB2AA42A8E2A772A602A492A322A1B2A0429ED29D729C029A9"
// synthesis attribute INIT_28 of requantizer_coefficient_RAM is "256'h2C712C5A2C432C2C2C152BFE2BE72BCF2BB82BA12B8A2B732B5C2B452B2E2B17"
// synthesis attribute INIT_29 of requantizer_coefficient_RAM is "256'h2DE52DCE2DB72D9F2D882D712D592D422D2B2D142CFC2CE52CCE2CB72CA02C88"
// synthesis attribute INIT_2A of requantizer_coefficient_RAM is "256'h2F5C2F452F2D2F162EFE2EE72ECF2EB82EA02E892E722E5A2E432E2B2E142DFD"
// synthesis attribute INIT_2B of requantizer_coefficient_RAM is "256'h30D630BF30A7308F3077306030483031301930012FEA2FD22FBB2FA32F8B2F74"
// synthesis attribute INIT_2C of requantizer_coefficient_RAM is "256'h3253323B3223320B31F431DC31C431AC3194317C3165314D3135311D310630EE"
// synthesis attribute INIT_2D of requantizer_coefficient_RAM is "256'h33D333BB33A3338B3373335B3343332B331332FB32E332CB32B3329B3283326B"
// synthesis attribute INIT_2E of requantizer_coefficient_RAM is "256'h3555353D3525350C34F434DC34C434AC3494347B3463344B3433341B340333EB"
// synthesis attribute INIT_2F of requantizer_coefficient_RAM is "256'h36DA36C236AA36913679366036483630361735FF35E735CE35B6359E3586356D"
// synthesis attribute INIT_30 of requantizer_coefficient_RAM is "256'h3862384A38313819380037E737CF37B6379E3785376D3755373C3724370B36F3"
// synthesis attribute INIT_31 of requantizer_coefficient_RAM is "256'h39ED39D439BB39A3398A3971395939403927390F38F638DD38C538AC3893387B"
// synthesis attribute INIT_32 of requantizer_coefficient_RAM is "256'h3B7A3B613B483B2F3B173AFE3AE53ACC3AB33A9A3A813A693A503A373A1E3A06"
// synthesis attribute INIT_33 of requantizer_coefficient_RAM is "256'h3D0A3CF13CD83CBF3CA63C8D3C743C5B3C423C293C103BF73BDE3BC53BAC3B93"
// synthesis attribute INIT_34 of requantizer_coefficient_RAM is "256'h3E9C3E833E6A3E513E373E1E3E053DEC3DD33DBA3DA13D873D6E3D553D3C3D23"
// synthesis attribute INIT_35 of requantizer_coefficient_RAM is "256'h2019200C3FFF3FE53FCC3FB23F993F803F663F4D3F343F1B3F013EE83ECF3EB6"
// synthesis attribute INIT_36 of requantizer_coefficient_RAM is "256'h20E520D820CB20BE20B220A52098208B207F207220652058204C203F20322026"
// synthesis attribute INIT_37 of requantizer_coefficient_RAM is "256'h21B221A52198218B217E217121652158214B213E213121252118210B20FE20F1"
// synthesis attribute INIT_38 of requantizer_coefficient_RAM is "256'h2280227322662259224C223F223222252219220C21FF21F221E521D821CB21BE"
// synthesis attribute INIT_39 of requantizer_coefficient_RAM is "256'h234F234223352328231B230E230122F422E722DA22CD22C022B422A7229A228D"
// synthesis attribute INIT_3A of requantizer_coefficient_RAM is "256'h24202413240623F923EC23DE23D123C423B723AA239D2390238323762369235C"
// synthesis attribute INIT_3B of requantizer_coefficient_RAM is "256'h24F224E424D724CA24BD24B024A324962489247B246E246124542447243A242D"
// synthesis attribute INIT_3C of requantizer_coefficient_RAM is "256'h25C525B725AA259D2590258325752568255B254E2541253325262519250C24FF"
// synthesis attribute INIT_3D of requantizer_coefficient_RAM is "256'h2699268B267E2671266426562649263C262E26212614260725F925EC25DF25D2"
// synthesis attribute INIT_3E of requantizer_coefficient_RAM is "256'h276E2761275327462739272B271E2710270326F626E926DB26CE26C126B326A6"
// synthesis attribute INIT_3F of requantizer_coefficient_RAM is "256'h284428372829281C280F280127F427E627D927CC27BE27B127A327962789277B"

// synthesis translate_off

defparam requantizer_coefficient_RAM.INIT_00 = 256'h24FF_21BE_3D23_36F3_30EE_2B17_2572_2000_3590_2B9D_2234_32CC_229E_2852_1000_0000;
defparam requantizer_coefficient_RAM.INIT_01 = 256'h30B1_2E9C_2C8D_2A84_2880_2684_248D_229E_20B5_3DA6_39F0_364A_32B4_2F2D_2BB7_2852;
defparam requantizer_coefficient_RAM.INIT_02 = 256'h2A68_2935_2804_26D6_25AA_2480_2359_2234_2111_3FE1_3DA6_3B70_393F_3713_34ED_32CC;
defparam requantizer_coefficient_RAM.INIT_03 = 256'h3EAC_3D59_3C09_3ABA_396C_3821_36D8_3590_344B_3307_31C6_3086_2F49_2E0D_2CD4_2B9D;
defparam requantizer_coefficient_RAM.INIT_04 = 256'h2A60_29A9_28F3_283E_278A_26D6_2623_2572_24C0_2410_2361_22B2_2204_2158_20AC_2000;
defparam requantizer_coefficient_RAM.INIT_05 = 256'h3630_356D_34AC_33EB_332B_326B_31AC_30EE_3031_2F74_2EB8_2DFD_2D42_2C88_2BCF_2B17;
defparam requantizer_coefficient_RAM.INIT_06 = 256'h2158_20F1_208B_2026_3F80_3EB6_3DEC_3D23_3C5B_3B93_3ACC_3A06_3940_387B_37B6_36F3;
defparam requantizer_coefficient_RAM.INIT_07 = 256'h27E6_277B_2710_26A6_263C_25D2_2568_24FF_2496_242D_23C4_235C_22F4_228D_2225_21BE;
defparam requantizer_coefficient_RAM.INIT_08 = 256'h2EBD_2E4E_2DDF_2D70_2D01_2C93_2C25_2BB7_2B49_2ADC_2A6F_2A02_2996_2929_28BD_2852;
defparam requantizer_coefficient_RAM.INIT_09 = 256'h35D7_3563_34F0_347D_340A_3398_3326_32B4_3242_31D0_315F_30EE_307D_300D_2F9D_2F2D;
defparam requantizer_coefficient_RAM.INIT_0A = 256'h3D2E_3CB7_3C40_3BC9_3B53_3ADC_3A66_39F0_397B_3906_3890_381B_37A7_3732_36BE_364A;
defparam requantizer_coefficient_RAM.INIT_0B = 256'h2260_2223_21E6_21A8_216B_212E_20F2_20B5_2078_203C_3FFE_3F86_3F0D_3E95_3E1D_3DA6;
defparam requantizer_coefficient_RAM.INIT_0C = 256'h2645_2605_25C7_2588_2549_250A_24CC_248D_244F_2411_23D3_2395_2357_2319_22DB_229E;
defparam requantizer_coefficient_RAM.INIT_0D = 256'h2A43_2A02_29C2_2981_2941_2901_28C1_2880_2841_2801_27C1_2781_2742_2702_26C3_2684;
defparam requantizer_coefficient_RAM.INIT_0E = 256'h2E5A_2E18_2DD6_2D94_2D52_2D10_2CCF_2C8D_2C4B_2C0A_2BC9_2B88_2B46_2B05_2AC4_2A84;
defparam requantizer_coefficient_RAM.INIT_0F = 256'h3289_3245_3202_31BE_317B_3138_30F5_30B1_306F_302C_2FE9_2FA6_2F64_2F21_2EDF_2E9C;
defparam requantizer_coefficient_RAM.INIT_10 = 256'h36CE_3689_3644_3600_35BB_3576_3532_34ED_34A9_3464_3420_33DC_3398_3354_3310_32CC;
defparam requantizer_coefficient_RAM.INIT_11 = 256'h3B29_3AE3_3A9D_3A57_3A11_39CB_3985_393F_38F9_38B3_386E_3828_37E3_379E_3758_3713;
defparam requantizer_coefficient_RAM.INIT_12 = 256'h3F99_3F52_3F0A_3EC3_3E7C_3E34_3DED_3DA6_3D5F_3D18_3CD1_3C8A_3C43_3BFD_3BB6_3B70;
defparam requantizer_coefficient_RAM.INIT_13 = 256'h220F_21EB_21C6_21A2_217E_2159_2135_2111_20ED_20C9_20A5_2081_205D_2039_2015_3FE1;
defparam requantizer_coefficient_RAM.INIT_14 = 256'h245B_2436_2411_23EC_23C7_23A2_237D_2359_2334_230F_22EA_22C6_22A1_227D_2258_2234;
defparam requantizer_coefficient_RAM.INIT_15 = 256'h26B0_268B_2665_2640_261A_25F5_25CF_25AA_2584_255F_253A_2515_24EF_24CA_24A5_2480;
defparam requantizer_coefficient_RAM.INIT_16 = 256'h290F_28E9_28C2_289C_2876_2850_282A_2804_27DE_27B9_2793_276D_2747_2721_26FC_26D6;
defparam requantizer_coefficient_RAM.INIT_17 = 256'h2B76_2B4F_2B29_2B02_2ADB_2AB5_2A8E_2A68_2A41_2A1B_29F5_29CE_29A8_2981_295B_2935;
defparam requantizer_coefficient_RAM.INIT_18 = 256'h2DE6_2DBF_2D98_2D70_2D49_2D22_2CFB_2CD4_2CAD_2C86_2C5F_2C38_2C11_2BEA_2BC4_2B9D;
defparam requantizer_coefficient_RAM.INIT_19 = 256'h305E_3037_300F_2FE7_2FC0_2F98_2F70_2F49_2F21_2EFA_2ED2_2EAB_2E83_2E5C_2E35_2E0D;
defparam requantizer_coefficient_RAM.INIT_1A = 256'h32DF_32B7_328F_3266_323E_3216_31EE_31C6_319E_3176_314E_3126_30FE_30D6_30AE_3086;
defparam requantizer_coefficient_RAM.INIT_1B = 256'h3568_353F_3516_34ED_34C5_349C_3473_344B_3422_33FA_33D1_33A9_3380_3358_3330_3307;
defparam requantizer_coefficient_RAM.INIT_1C = 256'h37F8_37CF_37A5_377C_3753_372A_3701_36D8_36AF_3686_365D_3634_360B_35E2_35B9_3590;
defparam requantizer_coefficient_RAM.INIT_1D = 256'h3A90_3A66_3A3C_3A13_39E9_39C0_3996_396C_3943_3919_38F0_38C7_389D_3874_384A_3821;
defparam requantizer_coefficient_RAM.INIT_1E = 256'h3D2F_3D05_3CDB_3CB1_3C87_3C5D_3C33_3C09_3BDF_3BB5_3B8B_3B61_3B37_3B0D_3AE3_3ABA;
defparam requantizer_coefficient_RAM.INIT_1F = 256'h3FD6_3FAB_3F81_3F56_3F2C_3F01_3ED7_3EAC_3E82_3E57_3E2D_3E03_3DD8_3DAE_3D84_3D59;
defparam requantizer_coefficient_RAM.INIT_20 = 256'h2142_212D_2117_2101_20EC_20D7_20C1_20AC_2096_2081_206B_2056_2041_202B_2016_2000;
defparam requantizer_coefficient_RAM.INIT_21 = 256'h229C_2287_2271_225B_2246_2230_221A_2204_21EF_21D9_21C4_21AE_2198_2183_216D_2158;
defparam requantizer_coefficient_RAM.INIT_22 = 256'h23FA_23E4_23CE_23B8_23A2_238D_2377_2361_234B_2335_231F_2309_22F4_22DE_22C8_22B2;
defparam requantizer_coefficient_RAM.INIT_23 = 256'h255B_2545_252F_2519_2503_24ED_24D7_24C0_24AA_2494_247E_2468_2452_243C_2426_2410;
defparam requantizer_coefficient_RAM.INIT_24 = 256'h26C0_26A9_2693_267D_2666_2650_263A_2623_260D_25F7_25E1_25CA_25B4_259E_2588_2572;
defparam requantizer_coefficient_RAM.INIT_25 = 256'h2827_2811_27FA_27E4_27CD_27B7_27A0_278A_2773_275D_2746_2730_2719_2703_26ED_26D6;
defparam requantizer_coefficient_RAM.INIT_26 = 256'h2992_297C_2965_294E_2937_2921_290A_28F3_28DC_28C6_28AF_2898_2882_286B_2855_283E;
defparam requantizer_coefficient_RAM.INIT_27 = 256'h2B00_2AE9_2AD2_2ABB_2AA4_2A8E_2A77_2A60_2A49_2A32_2A1B_2A04_29ED_29D7_29C0_29A9;
defparam requantizer_coefficient_RAM.INIT_28 = 256'h2C71_2C5A_2C43_2C2C_2C15_2BFE_2BE7_2BCF_2BB8_2BA1_2B8A_2B73_2B5C_2B45_2B2E_2B17;
defparam requantizer_coefficient_RAM.INIT_29 = 256'h2DE5_2DCE_2DB7_2D9F_2D88_2D71_2D59_2D42_2D2B_2D14_2CFC_2CE5_2CCE_2CB7_2CA0_2C88;
defparam requantizer_coefficient_RAM.INIT_2A = 256'h2F5C_2F45_2F2D_2F16_2EFE_2EE7_2ECF_2EB8_2EA0_2E89_2E72_2E5A_2E43_2E2B_2E14_2DFD;
defparam requantizer_coefficient_RAM.INIT_2B = 256'h30D6_30BF_30A7_308F_3077_3060_3048_3031_3019_3001_2FEA_2FD2_2FBB_2FA3_2F8B_2F74;
defparam requantizer_coefficient_RAM.INIT_2C = 256'h3253_323B_3223_320B_31F4_31DC_31C4_31AC_3194_317C_3165_314D_3135_311D_3106_30EE;
defparam requantizer_coefficient_RAM.INIT_2D = 256'h33D3_33BB_33A3_338B_3373_335B_3343_332B_3313_32FB_32E3_32CB_32B3_329B_3283_326B;
defparam requantizer_coefficient_RAM.INIT_2E = 256'h3555_353D_3525_350C_34F4_34DC_34C4_34AC_3494_347B_3463_344B_3433_341B_3403_33EB;
defparam requantizer_coefficient_RAM.INIT_2F = 256'h36DA_36C2_36AA_3691_3679_3660_3648_3630_3617_35FF_35E7_35CE_35B6_359E_3586_356D;
defparam requantizer_coefficient_RAM.INIT_30 = 256'h3862_384A_3831_3819_3800_37E7_37CF_37B6_379E_3785_376D_3755_373C_3724_370B_36F3;
defparam requantizer_coefficient_RAM.INIT_31 = 256'h39ED_39D4_39BB_39A3_398A_3971_3959_3940_3927_390F_38F6_38DD_38C5_38AC_3893_387B;
defparam requantizer_coefficient_RAM.INIT_32 = 256'h3B7A_3B61_3B48_3B2F_3B17_3AFE_3AE5_3ACC_3AB3_3A9A_3A81_3A69_3A50_3A37_3A1E_3A06;
defparam requantizer_coefficient_RAM.INIT_33 = 256'h3D0A_3CF1_3CD8_3CBF_3CA6_3C8D_3C74_3C5B_3C42_3C29_3C10_3BF7_3BDE_3BC5_3BAC_3B93;
defparam requantizer_coefficient_RAM.INIT_34 = 256'h3E9C_3E83_3E6A_3E51_3E37_3E1E_3E05_3DEC_3DD3_3DBA_3DA1_3D87_3D6E_3D55_3D3C_3D23;
defparam requantizer_coefficient_RAM.INIT_35 = 256'h2019_200C_3FFF_3FE5_3FCC_3FB2_3F99_3F80_3F66_3F4D_3F34_3F1B_3F01_3EE8_3ECF_3EB6;
defparam requantizer_coefficient_RAM.INIT_36 = 256'h20E5_20D8_20CB_20BE_20B2_20A5_2098_208B_207F_2072_2065_2058_204C_203F_2032_2026;
defparam requantizer_coefficient_RAM.INIT_37 = 256'h21B2_21A5_2198_218B_217E_2171_2165_2158_214B_213E_2131_2125_2118_210B_20FE_20F1;
defparam requantizer_coefficient_RAM.INIT_38 = 256'h2280_2273_2266_2259_224C_223F_2232_2225_2219_220C_21FF_21F2_21E5_21D8_21CB_21BE;
defparam requantizer_coefficient_RAM.INIT_39 = 256'h234F_2342_2335_2328_231B_230E_2301_22F4_22E7_22DA_22CD_22C0_22B4_22A7_229A_228D;
defparam requantizer_coefficient_RAM.INIT_3A = 256'h2420_2413_2406_23F9_23EC_23DE_23D1_23C4_23B7_23AA_239D_2390_2383_2376_2369_235C;
defparam requantizer_coefficient_RAM.INIT_3B = 256'h24F2_24E4_24D7_24CA_24BD_24B0_24A3_2496_2489_247B_246E_2461_2454_2447_243A_242D;
defparam requantizer_coefficient_RAM.INIT_3C = 256'h25C5_25B7_25AA_259D_2590_2583_2575_2568_255B_254E_2541_2533_2526_2519_250C_24FF;
defparam requantizer_coefficient_RAM.INIT_3D = 256'h2699_268B_267E_2671_2664_2656_2649_263C_262E_2621_2614_2607_25F9_25EC_25DF_25D2;
defparam requantizer_coefficient_RAM.INIT_3E = 256'h276E_2761_2753_2746_2739_272B_271E_2710_2703_26F6_26E9_26DB_26CE_26C1_26B3_26A6;
defparam requantizer_coefficient_RAM.INIT_3F = 256'h2844_2837_2829_281C_280F_2801_27F4_27E6_27D9_27CC_27BE_27B1_27A3_2796_2789_277B;

// synthesis translate_on

endmodule
